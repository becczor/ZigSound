--------------------------------------------------------------------------------
-- SOUND
-- Rebecca Lindblom
-- 31-mars-2017
-- Version 1.0


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type and various arithmetic operations

-- entity
entity SOUND is
port (
    clk                 : in std_logic;                      -- system clock (100 MHz)
    rst                 : in std_logic;                      -- reset signal
    goal_pos            : in signed(17 downto 0);  -- goal position
    curr_pos            : in signed(17 downto 0);  -- current position
    channel             : in std_logic;                      -- deciding which of the two sound that should be played, 0 = curr, 1 = goal.
    sound_data          : out std_logic);                    -- output to speaker
    --sound_enable        : in std_logic;                      -- possible for later to add on/off for sound
end SOUND;

-- architecture
architecture behavioral of SOUND is
    
    signal goal_x       : signed(5 downto 0);
    signal curr_x       : signed(5 downto 0);
   
    signal goal_y       : signed(4 downto 0);
    signal curr_y       : signed(4 downto 0);

    signal x            : signed(5 downto 0);         -- x-position for playing
    signal y            : signed(4 downto 0);         -- y-position for playing

    signal beat         : signed(19 downto 0);        -- Divided value for desired frequency for beat at position
    signal freq         : signed(10 downto 0);        -- Divided value for desired frequency for freq at position

    signal clk_div_beat : signed(19 downto 0);        -- Dividing clock for beat
    signal clk_div_freq : signed(10 downto 0);        -- Dividing clock for freq

    signal clk_beat     : std_logic;                            -- Clock signal for beat
    signal clk_freq     : std_logic;                            -- Clock signal for freq

    -- Flip flops
    signal q_beat       : std_logic := '0';                       -- Beat flip flop
    signal q_beat_plus  : std_logic := '0';    
    
    signal q_freq       : std_logic := '0';                       -- Freq flip flop
    signal q_freq_plus  : std_logic := '0';     

begin

    -- Set signals for playing sound
    process(clk)
    begin
        if rising_edge(clk) then
            if rst='1' then
                x <= "000000";
                y <= "00000";
            elsif channel = '1' then
                x <= goal_x;
                y <= goal_y;
            else
                x <= curr_x;
                y <= curr_y;
            end if;
        end if;
    end process;

    -- Transfer position data to internal signals
    process(clk)
    begin
        if rising_edge(clk) then
            -- Should look at registers all the time, even at reset
            goal_x <= goal_pos(14 downto 9);
            goal_y <= goal_pos(4 downto 0);
            curr_x <= curr_pos(14 downto 9);
            curr_y <= curr_pos(4 downto 0);
        end if;
    end process;


    -- y position -> beat value for toggle clk_beat
    -- follows beat = round(100000000 / (0.555764 * exp(0.0980482 * y)))
    -- See list of Hz-values in frequencies.txt
    -- Position is 0 at top of screen
    with y select
      beat <=
      1000000 when "11101",--29,
      789474  when "11100",--28,
      652174  when "11011",--27,
      555556  when "11010",--26,
      483871  when "11001",--25,
      428571  when "11000",--24,
      384615  when "10111",--23,
      348837  when "10110",--22,
      319149  when "10101",--21,
      294118  when "10100",--20,
      272727  when "10011",--19,
      250000  when "10010",--18,
      230769  when "10001",--17,
      214286  when "10000",--16,
      197368  when "01111",--15,
      180723  when "01110",--14,
      166667  when "01101",--13,
      153846  when "01100",--12,
      142180  when "01011",--11,
      130435  when "01010",--10,
      119048  when "01001",--9,
      109091  when "01000",--8,
      100000  when "00111",--7,
      90909   when "00110"--6,
      81081   when "00101",--5,
      73171   when "00100",--4,
      65217   when "00011",--3,
      57692   when "00010",--2,
      50847   when "00001",--1,
      45455   when "00000",--0,
      1       when others;

    -- x-position -> freq value for toggle clk_freq
    -- Follows freq <= round(100000000/ (300 + 25*x)
    -- See list of Hz-values in frequencies.txt
    -- Position is 0 at left of screen
    with x select
      freq <=
      1538 when "000000",--0,
      1429 when "000001",--1,
      1333 when "000010",--2,
      1250 when "000011",--3,
      1176 when "000100",--4,
      1111 when "000101",--5,
      1053 when "000110",--6,
      1000 when "000111",--7,
      952  when "001000",--8,
      909  when "001001",--9,
      870  when "001010",--10,
      833  when "001011",--11,
      800  when "001100",--12,
      769  when "001101",--13,
      741  when "001110",--14,
      714  when "001111",--15,
      690  when "010000",--16,
      667  when "010001",--17,
      645  when "010010",--18,
      625  when "010011",--19,
      606  when "010100",--20,
      588  when "010101",--21,
      571  when "010110",--22,
      556  when "010111",--23,
      541  when "011000",--24,
      526  when "011001",--25,
      513  when "011010",--26,
      500  when "011011",--27,
      488  when "011100",--28
      476  when "011101",--29,
      465  when "011110",--30,
      455  when "011111",--31,
      444  when "100000",--32,
      435  when "100001",--33,
      426  when "100010",--34,
      417  when "100011",--35,
      408  when "100100",--36,
      400  when "100101",--37,
      392  when "100110",--38,
      385  when "100111",--39,
      1    when others;

        
    -- Clock divisor
    -- Divide system clock (100 MHz) by beat and freq
    process(clk) begin
        if rising_edge(clk) then
            if rst='1' then
                clk_div_beat <= (others => '0');
                clk_div_freq <= (others => '0');
            elsif clk_div_beat = beat then
                clk_div_beat <= 0;
            elsif clk_div_freq = beat then
                clk_div_freq <= 0;
            else
                clk_div_beat <= clk_div_beat + 1;
                clk_div_freq <= clk_div_freq + 1;
            end if;
        end if;
    end process;

    -- Toggle sound clocks to get 50% duty cycle
    clk_beat <= not clk_beat when (clk_beat_div < beat) else clk_beat;
    clk_freq <= not clk_freq when (clk_freq_div < freq) else clk_freq;


    -- Beat flip flop
    process(clk_beat) begin
        if rising_edge(clk_beat) then
            if rst='1' then
                q_beat <= 0;
            else
                q_beat <= q_beat_plus;
            end if;
        end if;
    end process;

    -- Freq flip flop
    process(clk_freq) begin
        if rising_edge(clk_beat) then
            if rst='1' then
                q_freq <= 0;
            else
                q_freq <= q_freq_plus;
            end if;
        end if;
    end process;
        
    --q_beat_plus <= sound_enable and not q_beat;
    q_beat_plus <= not q_beat;
    q_freq_plus <= q_beat and not q_freq;
  
end behavioral;
