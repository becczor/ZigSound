sabse455@mux2-09.edu.isy.liu.se.5489:1493300119