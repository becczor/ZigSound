library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

--*****************
--* CPU interface *
--*****************
entity CPU is
    port(
        clk                 : in std_logic;
        rst                 : in std_logic;
        uAddr               : out unsigned(6 downto 0);
        uData               : in unsigned(24 downto 0);
        pAddr               : out signed(7 downto 0);
        pData               : in signed(17 downto 0);
        PS2cmd              : in unsigned(17 downto 0);
		move_req_out        : out std_logic;
		upd_sound_icon_out  : out std_logic;
		move_resp           : in std_logic;
		curr_pos_out        : out signed(17 downto 0);
		next_pos_out        : out signed(17 downto 0);
        goal_pos_out        : out signed(17 downto 0);
		sel_track_out       : out unsigned(1 downto 0);
		sel_sound_out       : out std_logic;
		goal_reached_out    : out std_logic;
		showing_goal_msg    : in std_logic;
		disp_goal_pos_out   : out std_logic;
        score_out           : out unsigned(5 downto 0)
        );
end CPU;

architecture Behavioral of CPU is

    --****************
    --* Port aliases *
    --****************
    alias uM                : unsigned(24 downto 0) is uData(24 downto 0);
    alias PM                : signed(17 downto 0) is pData(17 downto 0);
    
    --*****************************
    --* Micro Instruction Aliases *
    --*****************************
    alias ALU               : unsigned(3 downto 0) is uM(24 downto 21);  -- ALU    
    alias TB                : unsigned(2 downto 0) is uM(20 downto 18);  -- To bus
    alias FB                : unsigned(2 downto 0) is uM(17 downto 15);  -- From bus
    alias S                 : std_logic is uM(14);                       -- S-bit
    alias P                 : std_logic is uM(13);                       -- P-bit
    alias LC                : unsigned(1 downto 0) is uM(12 downto 11);  -- LC
    alias SEQ               : unsigned(3 downto 0) is uM(10 downto 7);   -- SEQ
    alias MICROADDR         : unsigned(6 downto 0) is uM(6 downto 0);    -- Micro address
    
    --**************************************
    --* Program Memory Instruction Signals *
    --**************************************
    signal OP               : signed(4 downto 0);  -- Operation    
    signal GRX              : signed(2 downto 0);  -- Register    
    signal M                : signed(1 downto 0);  -- Addressing mode        
    signal ADDR             : signed(7 downto 0);  -- Address field    
	
    --****************
    --* Flag Signals *
    --****************
	signal flag_Z           : std_logic := '0';  -- Zero
	signal flag_N           : std_logic := '0';  -- Negative
	signal flag_C           : std_logic := '0';  -- NOT ALWAYS BEING DETECTED ATM
	signal flag_O           : std_logic := '0';  -- NOT BEING DETECTED ATM
	signal flag_L           : std_logic := '0';  -- 1 if LC_cnt = 0 (done)
    signal flag_G           : std_logic := '0';  -- Goal reached
    signal flag_S           : std_logic := '0';  -- VGA_MOTOR is showing goal message

    --****************************
    --* Outgoing signals signals *
    --****************************
    -- To GPU
    signal MOVE_REQ         : std_logic := '0';  -- Move request (move_req_out)
    signal UPD_SOUND_ICON   : std_logic := '0';  -- Signal for updating sound icon
    signal CURR_POS         : signed(17 downto 0) := "000000001000000001"; -- Current Position (curr_pos_out)
    signal NEXT_POS         : signed(17 downto 0) := "000000001000000001";  -- Next Postition (next_pos_out)
    signal SEL_TRACK        : signed(1 downto 0) := "00";  -- Track select (sel_track_out)
    -- To SOUND
    signal SEL_SOUND        : std_logic := '0'; -- Sound select (sel_sound_out)
    signal DISP_GOAL_POS    : std_logic := '0'; -- Display goal pos on screen (disp_goal_pos_out)
    signal GOAL_POS         : signed(17 downto 0) := (others => '0');  -- Goal position (goal_pos_out)
    signal RND_GOAL_POS     : signed(17 downto 0) := (others => '0');
    signal SCORE            : signed(17 downto 0) := (others => '0');
    signal WON              : std_logic := '0'; -- LSB signals that goal_pos was found

    --***************
    --* CPU Signals *
    --***************
    signal PC               : signed(7 downto 0) := (others => '0'); -- Program Counter
    signal uPC              : unsigned(6 downto 0) := (others => '0'); -- Micro Program Counter (uAddr)
	signal IR               : signed(17 downto 0) := (others => '0'); -- Instruction Register 
	signal DATA_BUS         : signed(17 downto 0) := (others => '0'); -- Data Bus
    signal ASR              : signed(7 downto 0) := (others => '0');  -- (pAddr)
    signal AR               : signed(17 downto 0) := (others => '0');
    signal GR0              : signed(17 downto 0) := (others => '0');
    signal GR1              : signed(17 downto 0) := (others => '0');
    signal GR2              : signed(17 downto 0) := (others => '0');
    signal GR3              : signed(17 downto 0) := (others => '0');
    signal NEXT_TRACK       : signed(17 downto 0) := (others => '1');
    
    --******************
    --* Signal aliases *
    --******************
    alias CURR_XPOS         : signed(5 downto 0) is CURR_POS(14 downto 9);
    alias CURR_YPOS         : signed(4 downto 0) is CURR_POS(4 downto 0);
    alias NEXT_XPOS         : signed(5 downto 0) is NEXT_POS(14 downto 9);
    alias NEXT_YPOS         : signed(4 downto 0) is NEXT_POS(4 downto 0);
    alias GOAL_XPOS         : signed(5 downto 0) is GOAL_POS(14 downto 9);
    alias GOAL_YPOS         : signed(4 downto 0) is GOAL_POS(4 downto 0);
    alias key_code          : unsigned(2 downto 0) is PS2cmd(2 downto 0);

    --************
    --* Counters *
    --************
    signal free_pos_lmt     : signed(10 downto 0) := (others => '0');
    signal free_pos_cnt     : signed(10 downto 0) := (others => '0');
    signal dly_cnt          : unsigned(2 downto 0) := (others => '0');
    signal LC_cnt           : signed(16 downto 0) := (others => '0');

     --TEST                             
    --signal test_led_counter             : unsigned(25 downto 0);
    --signal test_signal                  : std_logic;
    --signal working                      : std_logic;

    --****************************************************************************
	--* uAddr_instr : Array of uAddresses where each instruction begins in uMem. *
	--****************************************************************************
	type uAddr_instr_t is array (0 to 31) of unsigned(6 downto 0);
	constant uAddr_instr_c : uAddr_instr_t := 
	-- OP consists of 5 bits, so the maximum amount of instructions is 32.
    -------- µStartAddr ------- µInstr ----------- OP ---
        ("0001010",--x"0A", -- LOAD             "00000" 0
         "0001011",--x"0B", -- STORE            "00001" 1
         "0001100",--x"0C", -- ADD              "00010" 2
         "0001111",--x"0F", -- SUB              "00011" 3
         "0010010",--x"12", -- AND              "00100" 4
         "0010101",--x"15", -- LSR              "00101" 5
         "0011011",--x"1B", -- BRA              "00110" 6
         "0011110",--x"1E", -- CMP              "00111" 7
         "0100000",--x"20", -- BNE              "01000" 8
         "0100010",--x"22", -- BGT              "01001" 9
         "0101001",--x"29", -- BGE              "01010" 10
         "0101110",--x"2E", -- HALT             "01011" 11
         "0101111",--x"2F", -- BCT              "01100" 12
         "0110001",--x"31", -- SETRNDGOALPOS    "01101" 13 --GRX MUST BE "100"!
         "0110010",--x"32", -- SHOWGOALMSG      "01110" 14
         "0110100",--x"34", -- HIDEGOALMSG      "01111" 15
         "0110110",--x"36", -- WAIT             "10000" 16
         "0111010",--x"3A", -- INCRSCORE        "10001" 17
         "0111101",--x"3D", -- SENDWONSIG       "10010" 18
         "1000001",--x"41", -- BSW              "10011" 19
         "1000011",--x"43", -- INCRTRACK        "10100" 20 --GRX MUST BE "101"!
         "0000000",--x"00", -- NULL             "10101" 21
         "0000000",--x"00", -- NULL             "10110" 22
         "0000000",--x"00", -- NULL             "10111" 23
         "0000000",--x"00", -- NULL             "11000" 24
         "0000000",--x"00", -- NULL             "11001" 25
         "0000000",--x"00", -- NULL             "11010" 26
         "0000000",--x"00", -- NULL             "11011" 27
         "0000000",--x"00", -- NULL             "11100" 28
         "0000000",--x"00", -- NULL             "11101" 29
         "0000000",--x"00", -- NULL             "11110" 30
         "0000000" --x"00"  -- NULL             "11111" 31
        );
    signal uAddr_instr : uAddr_instr_t := uAddr_instr_c;
    
    --**************************
    --* p_mem : Program Memory *
    --**************************
    type track_1_free_pos_mem_t is array (0 to 913) of signed(17 downto 0);
    constant track_1_free_pos_mem_c : track_1_free_pos_mem_t := (
        -- Row: 0
        -- Row: 1
        b"000000010000000001",b"000000011000000001",b"000000100000000001",b"000000101000000001",
        b"000000110000000001",b"000000111000000001",b"000001000000000001",b"000001001000000001",
        b"000001010000000001",b"000001011000000001",b"000001100000000001",b"000001101000000001",
        b"000001110000000001",b"000001111000000001",b"000010000000000001",b"000010001000000001",
        b"000010011000000001",b"000010100000000001",b"000010101000000001",b"000010110000000001",
        b"000011000000000001",b"000011001000000001",b"000011010000000001",b"000011011000000001",
        b"000011100000000001",b"000011101000000001",b"000011110000000001",b"000011111000000001",
        b"000100000000000001",b"000100001000000001",b"000100010000000001",b"000100011000000001",
        b"000100100000000001",b"000100101000000001",b"000100110000000001",
        -- Row: 2
        b"000000001000000010",b"000000010000000010",b"000000011000000010",b"000000100000000010",
        b"000000101000000010",b"000000110000000010",b"000000111000000010",b"000001000000000010",
        b"000001001000000010",b"000001010000000010",b"000001011000000010",b"000001100000000010",
        b"000001101000000010",b"000001110000000010",b"000010000000000010",b"000010001000000010",
        b"000010010000000010",b"000010011000000010",b"000010100000000010",b"000010101000000010",
        b"000010111000000010",b"000011000000000010",b"000011001000000010",b"000011010000000010",
        b"000011011000000010",b"000011101000000010",b"000011110000000010",b"000011111000000010",
        b"000100000000000010",b"000100001000000010",b"000100010000000010",b"000100011000000010",
        b"000100100000000010",b"000100101000000010",
        -- Row: 3
        b"000000001000000011",b"000000010000000011",b"000000011000000011",b"000000100000000011",
        b"000000101000000011",b"000000111000000011",b"000001000000000011",b"000001001000000011",
        b"000001011000000011",b"000001100000000011",b"000001101000000011",b"000001110000000011",
        b"000001111000000011",b"000010001000000011",b"000010010000000011",b"000010011000000011",
        b"000010100000000011",b"000010101000000011",b"000010110000000011",b"000010111000000011",
        b"000011000000000011",b"000011001000000011",b"000011010000000011",b"000011100000000011",
        b"000011101000000011",b"000011110000000011",b"000011111000000011",b"000100000000000011",
        b"000100010000000011",b"000100011000000011",b"000100110000000011",
        -- Row: 4
        b"000000001000000100",b"000000010000000100",b"000000011000000100",b"000000100000000100",
        b"000000101000000100",b"000000110000000100",b"000000111000000100",b"000001000000000100",
        b"000001001000000100",b"000001011000000100",b"000001100000000100",b"000001101000000100",
        b"000001110000000100",b"000001111000000100",b"000010000000000100",b"000010001000000100",
        b"000010010000000100",b"000010011000000100",b"000010100000000100",b"000010101000000100",
        b"000010110000000100",b"000010111000000100",b"000011001000000100",b"000011010000000100",
        b"000011011000000100",b"000011100000000100",b"000011101000000100",b"000011110000000100",
        b"000011111000000100",b"000100000000000100",b"000100001000000100",b"000100010000000100",
        b"000100011000000100",b"000100100000000100",b"000100101000000100",b"000100110000000100",
        -- Row: 5
        b"000000001000000101",b"000000011000000101",b"000000100000000101",b"000000101000000101",
        b"000000110000000101",b"000000111000000101",b"000001000000000101",b"000001001000000101",
        b"000001010000000101",b"000001011000000101",b"000001100000000101",b"000001101000000101",
        b"000001110000000101",b"000001111000000101",b"000010000000000101",b"000010001000000101",
        b"000010010000000101",b"000010011000000101",b"000010101000000101",b"000010110000000101",
        b"000011000000000101",b"000011001000000101",b"000011010000000101",b"000011011000000101",
        b"000011100000000101",b"000011101000000101",b"000011110000000101",b"000011111000000101",
        b"000100001000000101",b"000100010000000101",b"000100011000000101",b"000100100000000101",
        b"000100101000000101",b"000100110000000101",
        -- Row: 6
        b"000000001000000110",b"000000010000000110",b"000000101000000110",b"000000110000000110",
        b"000000111000000110",b"000001000000000110",b"000001001000000110",b"000001010000000110",
        b"000001011000000110",b"000001101000000110",b"000001110000000110",b"000001111000000110",
        b"000010000000000110",b"000010001000000110",b"000010010000000110",b"000010011000000110",
        b"000010100000000110",b"000010110000000110",b"000010111000000110",b"000011000000000110",
        b"000011001000000110",b"000011011000000110",b"000011100000000110",b"000011101000000110",
        b"000011110000000110",b"000100000000000110",b"000100001000000110",b"000100010000000110",
        b"000100011000000110",b"000100101000000110",b"000100110000000110",
        -- Row: 7
        b"000000001000000111",b"000000010000000111",b"000000100000000111",b"000000101000000111",
        b"000000110000000111",b"000000111000000111",b"000001000000000111",b"000001001000000111",
        b"000001010000000111",b"000001011000000111",b"000001100000000111",b"000001101000000111",
        b"000001110000000111",b"000001111000000111",b"000010001000000111",b"000010010000000111",
        b"000010011000000111",b"000010100000000111",b"000010101000000111",b"000010110000000111",
        b"000010111000000111",b"000011000000000111",b"000011001000000111",b"000011011000000111",
        b"000011100000000111",b"000011101000000111",b"000100000000000111",b"000100001000000111",
        b"000100010000000111",b"000100011000000111",b"000100100000000111",b"000100110000000111",
        -- Row: 8
        b"000000010000001000",b"000000011000001000",b"000000100000001000",b"000000101000001000",
        b"000000110000001000",b"000001000000001000",b"000001001000001000",b"000001010000001000",
        b"000001011000001000",b"000001100000001000",b"000001101000001000",b"000001110000001000",
        b"000010001000001000",b"000010010000001000",b"000010011000001000",b"000010100000001000",
        b"000010101000001000",b"000010110000001000",b"000010111000001000",b"000011000000001000",
        b"000011010000001000",b"000011011000001000",b"000011100000001000",b"000011101000001000",
        b"000011110000001000",b"000011111000001000",b"000100000000001000",b"000100001000001000",
        b"000100010000001000",b"000100011000001000",b"000100100000001000",b"000100101000001000",
        b"000100110000001000",
        -- Row: 9
        b"000000001000001001",b"000000010000001001",b"000000011000001001",b"000000100000001001",
        b"000000101000001001",b"000000110000001001",b"000000111000001001",b"000001001000001001",
        b"000001011000001001",b"000001100000001001",b"000001101000001001",b"000001110000001001",
        b"000001111000001001",b"000010000000001001",b"000010001000001001",b"000010010000001001",
        b"000010011000001001",b"000010100000001001",b"000010111000001001",b"000011000000001001",
        b"000011001000001001",b"000011010000001001",b"000011011000001001",b"000011100000001001",
        b"000011101000001001",b"000011110000001001",b"000011111000001001",b"000100000000001001",
        b"000100011000001001",b"000100100000001001",b"000100101000001001",b"000100110000001001",
        -- Row: 10
        b"000000001000001010",b"000000010000001010",b"000000011000001010",b"000000100000001010",
        b"000000101000001010",b"000000110000001010",b"000001000000001010",b"000001011000001010",
        b"000001100000001010",b"000001101000001010",b"000001110000001010",b"000001111000001010",
        b"000010000000001010",b"000010001000001010",b"000010010000001010",b"000010011000001010",
        b"000010100000001010",b"000010101000001010",b"000011000000001010",b"000011001000001010",
        b"000011010000001010",b"000011011000001010",b"000011100000001010",b"000011111000001010",
        b"000100000000001010",b"000100001000001010",b"000100010000001010",b"000100011000001010",
        b"000100100000001010",b"000100101000001010",b"000100110000001010",
        -- Row: 11
        b"000000001000001011",b"000000011000001011",b"000000100000001011",b"000000101000001011",
        b"000000110000001011",b"000000111000001011",b"000001000000001011",b"000001010000001011",
        b"000001011000001011",b"000001100000001011",b"000001110000001011",b"000001111000001011",
        b"000010000000001011",b"000010001000001011",b"000010010000001011",b"000010100000001011",
        b"000010101000001011",b"000010110000001011",b"000010111000001011",b"000011000000001011",
        b"000011001000001011",b"000011010000001011",b"000011011000001011",b"000011100000001011",
        b"000011101000001011",b"000011110000001011",b"000011111000001011",b"000100000000001011",
        b"000100001000001011",b"000100010000001011",b"000100011000001011",b"000100100000001011",
        b"000100110000001011",
        -- Row: 12
        b"000000001000001100",b"000000010000001100",b"000000011000001100",b"000000100000001100",
        b"000000110000001100",b"000000111000001100",b"000001000000001100",b"000001001000001100",
        b"000001010000001100",b"000001011000001100",b"000001110000001100",b"000001111000001100",
        b"000010001000001100",b"000010010000001100",b"000010011000001100",b"000010101000001100",
        b"000010110000001100",b"000010111000001100",b"000011000000001100",b"000011001000001100",
        b"000011010000001100",b"000011100000001100",b"000011101000001100",b"000011110000001100",
        b"000011111000001100",b"000100001000001100",b"000100010000001100",b"000100011000001100",
        b"000100100000001100",b"000100101000001100",b"000100110000001100",
        -- Row: 13
        b"000000001000001101",b"000000010000001101",b"000000011000001101",b"000000100000001101",
        b"000000101000001101",b"000000110000001101",b"000000111000001101",b"000001000000001101",
        b"000001001000001101",b"000001010000001101",b"000001011000001101",b"000001100000001101",
        b"000001101000001101",b"000001110000001101",b"000001111000001101",b"000010000000001101",
        b"000010010000001101",b"000010011000001101",b"000010100000001101",b"000010110000001101",
        b"000010111000001101",b"000011000000001101",b"000011001000001101",b"000011011000001101",
        b"000011100000001101",b"000011101000001101",b"000011110000001101",b"000011111000001101",
        b"000100000000001101",b"000100001000001101",b"000100010000001101",b"000100100000001101",
        b"000100101000001101",b"000100110000001101",
        -- Row: 14
        b"000000001000001110",b"000000010000001110",b"000000011000001110",b"000000100000001110",
        b"000000101000001110",b"000000110000001110",b"000000111000001110",b"000001000000001110",
        b"000001001000001110",b"000001010000001110",b"000001011000001110",b"000001100000001110",
        b"000001101000001110",b"000001110000001110",b"000001111000001110",b"000010010000001110",
        b"000010011000001110",b"000010100000001110",b"000010101000001110",b"000010110000001110",
        b"000010111000001110",b"000011000000001110",b"000011001000001110",b"000011010000001110",
        b"000011011000001110",b"000011100000001110",b"000011101000001110",b"000011110000001110",
        b"000011111000001110",b"000100000000001110",b"000100001000001110",b"000100010000001110",
        b"000100011000001110",b"000100110000001110",
        -- Row: 15
        b"000000001000001111",b"000000010000001111",b"000000011000001111",b"000000101000001111",
        b"000000111000001111",b"000001000000001111",b"000001001000001111",b"000001010000001111",
        b"000001100000001111",b"000001101000001111",b"000001110000001111",b"000010000000001111",
        b"000010001000001111",b"000010010000001111",b"000010011000001111",b"000010100000001111",
        b"000010101000001111",b"000010110000001111",b"000011000000001111",b"000011001000001111",
        b"000011010000001111",b"000011011000001111",b"000011101000001111",b"000011110000001111",
        b"000100000000001111",b"000100001000001111",b"000100010000001111",b"000100011000001111",
        b"000100100000001111",b"000100101000001111",b"000100110000001111",
        -- Row: 16
        b"000000001000010000",b"000000010000010000",b"000000011000010000",b"000000100000010000",
        b"000000110000010000",b"000000111000010000",b"000001000000010000",b"000001011000010000",
        b"000001100000010000",b"000001101000010000",b"000001110000010000",b"000001111000010000",
        b"000010000000010000",b"000010001000010000",b"000010010000010000",b"000010011000010000",
        b"000010100000010000",b"000010101000010000",b"000010111000010000",b"000011000000010000",
        b"000011001000010000",b"000011010000010000",b"000011011000010000",b"000011100000010000",
        b"000011101000010000",b"000011110000010000",b"000100010000010000",b"000100011000010000",
        b"000100100000010000",b"000100101000010000",b"000100110000010000",
        -- Row: 17
        b"000000001000010001",b"000000011000010001",b"000000100000010001",b"000000101000010001",
        b"000000110000010001",b"000000111000010001",b"000001000000010001",b"000001001000010001",
        b"000001010000010001",b"000001100000010001",b"000001101000010001",b"000001110000010001",
        b"000001111000010001",b"000010000000010001",b"000010001000010001",b"000010010000010001",
        b"000010100000010001",b"000010101000010001",b"000010111000010001",b"000011000000010001",
        b"000011001000010001",b"000011010000010001",b"000011011000010001",b"000011100000010001",
        b"000011101000010001",b"000011110000010001",b"000011111000010001",b"000100000000010001",
        b"000100001000010001",b"000100010000010001",b"000100011000010001",b"000100100000010001",
        b"000100101000010001",
        -- Row: 18
        b"000000001000010010",b"000000010000010010",b"000000011000010010",b"000000100000010010",
        b"000000101000010010",b"000000110000010010",b"000000111000010010",b"000001000000010010",
        b"000001001000010010",b"000001010000010010",b"000001011000010010",b"000001100000010010",
        b"000001101000010010",b"000001110000010010",b"000001111000010010",b"000010000000010010",
        b"000010001000010010",b"000010011000010010",b"000010100000010010",b"000010101000010010",
        b"000010110000010010",b"000010111000010010",b"000011000000010010",b"000011001000010010",
        b"000011100000010010",b"000011101000010010",b"000011110000010010",b"000011111000010010",
        b"000100000000010010",b"000100001000010010",b"000100011000010010",b"000100100000010010",
        b"000100101000010010",b"000100110000010010",
        -- Row: 19
        b"000000001000010011",b"000000010000010011",b"000000011000010011",b"000000100000010011",
        b"000000101000010011",b"000000110000010011",b"000000111000010011",b"000001000000010011",
        b"000001001000010011",b"000001010000010011",b"000001011000010011",b"000001100000010011",
        b"000001101000010011",b"000001110000010011",b"000001111000010011",b"000010000000010011",
        b"000010001000010011",b"000010010000010011",b"000010100000010011",b"000010101000010011",
        b"000010110000010011",b"000010111000010011",b"000011000000010011",b"000011001000010011",
        b"000011010000010011",b"000011100000010011",b"000011101000010011",b"000011110000010011",
        b"000011111000010011",b"000100000000010011",b"000100010000010011",b"000100011000010011",
        b"000100100000010011",b"000100101000010011",b"000100110000010011",
        -- Row: 20
        b"000000001000010100",b"000000010000010100",b"000000011000010100",b"000000100000010100",
        b"000000111000010100",b"000001000000010100",b"000001001000010100",b"000001011000010100",
        b"000001100000010100",b"000001101000010100",b"000001110000010100",b"000010000000010100",
        b"000010001000010100",b"000010010000010100",b"000010011000010100",b"000010100000010100",
        b"000010101000010100",b"000010110000010100",b"000010111000010100",b"000011000000010100",
        b"000011001000010100",b"000011010000010100",b"000011011000010100",b"000011100000010100",
        b"000011101000010100",b"000011110000010100",b"000011111000010100",b"000100000000010100",
        b"000100001000010100",b"000100010000010100",b"000100011000010100",b"000100110000010100",
        -- Row: 21
        b"000000001000010101",b"000000010000010101",b"000000011000010101",b"000000110000010101",
        b"000000111000010101",b"000001000000010101",b"000001001000010101",b"000001010000010101",
        b"000001100000010101",b"000001101000010101",b"000001110000010101",b"000001111000010101",
        b"000010000000010101",b"000010001000010101",b"000010010000010101",b"000010011000010101",
        b"000010100000010101",b"000010101000010101",b"000010110000010101",b"000010111000010101",
        b"000011000000010101",b"000011001000010101",b"000011011000010101",b"000011100000010101",
        b"000011101000010101",b"000011111000010101",b"000100000000010101",b"000100001000010101",
        b"000100010000010101",b"000100011000010101",b"000100101000010101",b"000100110000010101",
        -- Row: 22
        b"000000001000010110",b"000000010000010110",b"000000100000010110",b"000000101000010110",
        b"000000110000010110",b"000000111000010110",b"000001000000010110",b"000001001000010110",
        b"000001010000010110",b"000001100000010110",b"000001101000010110",b"000001110000010110",
        b"000001111000010110",b"000010000000010110",b"000010001000010110",b"000010010000010110",
        b"000010011000010110",b"000010100000010110",b"000010110000010110",b"000010111000010110",
        b"000011001000010110",b"000011010000010110",b"000011011000010110",b"000011100000010110",
        b"000011101000010110",b"000011110000010110",b"000100000000010110",b"000100001000010110",
        b"000100010000010110",b"000100011000010110",b"000100100000010110",b"000100101000010110",
        b"000100110000010110",
        -- Row: 23
        b"000000001000010111",b"000000010000010111",b"000000100000010111",b"000000101000010111",
        b"000000110000010111",b"000000111000010111",b"000001000000010111",b"000001001000010111",
        b"000001010000010111",b"000001011000010111",b"000001100000010111",b"000001101000010111",
        b"000001110000010111",b"000010000000010111",b"000010001000010111",b"000010011000010111",
        b"000010100000010111",b"000010101000010111",b"000010110000010111",b"000011000000010111",
        b"000011001000010111",b"000011010000010111",b"000011011000010111",b"000011100000010111",
        b"000011101000010111",b"000011110000010111",b"000011111000010111",b"000100000000010111",
        b"000100001000010111",b"000100010000010111",b"000100011000010111",b"000100100000010111",
        b"000100101000010111",b"000100110000010111",
        -- Row: 24
        b"000000001000011000",b"000000100000011000",b"000000101000011000",b"000000111000011000",
        b"000001000000011000",b"000001001000011000",b"000001010000011000",b"000001011000011000",
        b"000001100000011000",b"000001101000011000",b"000001111000011000",b"000010000000011000",
        b"000010001000011000",b"000010011000011000",b"000010100000011000",b"000010101000011000",
        b"000010110000011000",b"000010111000011000",b"000011001000011000",b"000011010000011000",
        b"000011011000011000",b"000011101000011000",b"000011110000011000",b"000011111000011000",
        b"000100000000011000",b"000100010000011000",b"000100011000011000",b"000100101000011000",
        b"000100110000011000",
        -- Row: 25
        b"000000001000011001",b"000000010000011001",b"000000011000011001",b"000000100000011001",
        b"000000101000011001",b"000000110000011001",b"000000111000011001",b"000001000000011001",
        b"000001010000011001",b"000001011000011001",b"000001100000011001",b"000001101000011001",
        b"000001110000011001",b"000001111000011001",b"000010000000011001",b"000010001000011001",
        b"000010010000011001",b"000010100000011001",b"000010101000011001",b"000010110000011001",
        b"000010111000011001",b"000011000000011001",b"000011001000011001",b"000011010000011001",
        b"000011011000011001",b"000011101000011001",b"000011110000011001",b"000011111000011001",
        b"000100000000011001",b"000100001000011001",b"000100010000011001",b"000100011000011001",
        b"000100100000011001",b"000100110000011001",
        -- Row: 26
        b"000000001000011010",b"000000010000011010",b"000000011000011010",b"000000100000011010",
        b"000000101000011010",b"000000110000011010",b"000000111000011010",b"000001000000011010",
        b"000001001000011010",b"000001010000011010",b"000001011000011010",b"000001100000011010",
        b"000001101000011010",b"000001110000011010",b"000001111000011010",b"000010000000011010",
        b"000010001000011010",b"000010010000011010",b"000010100000011010",b"000010101000011010",
        b"000010110000011010",b"000010111000011010",b"000011000000011010",b"000011001000011010",
        b"000011010000011010",b"000011011000011010",b"000011100000011010",b"000011110000011010",
        b"000011111000011010",b"000100000000011010",b"000100001000011010",b"000100011000011010",
        b"000100100000011010",b"000100101000011010",b"000100110000011010",
        -- Row: 27
        b"000000001000011011",b"000000010000011011",b"000000011000011011",b"000000100000011011",
        b"000000111000011011",b"000001000000011011",b"000001001000011011",b"000001011000011011",
        b"000001100000011011",b"000001110000011011",b"000001111000011011",b"000010000000011011",
        b"000010001000011011",b"000010010000011011",b"000010011000011011",b"000010100000011011",
        b"000010101000011011",b"000010111000011011",b"000011000000011011",b"000011001000011011",
        b"000011011000011011",b"000011100000011011",b"000011101000011011",b"000011110000011011",
        b"000011111000011011",b"000100000000011011",b"000100001000011011",b"000100010000011011",
        b"000100100000011011",b"000100101000011011",
        -- Row: 28
        b"000000001000011100",b"000000011000011100",b"000000100000011100",b"000000101000011100",
        b"000000110000011100",b"000000111000011100",b"000001000000011100",b"000001010000011100",
        b"000001011000011100",b"000001100000011100",b"000001101000011100",b"000001111000011100",
        b"000010000000011100",b"000010010000011100",b"000010011000011100",b"000010100000011100",
        b"000010110000011100",b"000010111000011100",b"000011000000011100",b"000011001000011100",
        b"000011010000011100",b"000011100000011100",b"000011101000011100",b"000011110000011100",
        b"000011111000011100",b"000100001000011100",b"000100010000011100",b"000100011000011100",
        b"000100100000011100",b"000100101000011100"
        -- Row: 29
   
	        );
	
	    type track_2_free_pos_mem_t is array (0 to 886) of signed(17 downto 0);
	    constant track_2_free_pos_mem_c : track_2_free_pos_mem_t := (
           -- Row: 0
        -- Row: 1
        b"000000010000000001",b"000000011000000001",b"000000100000000001",b"000000101000000001",
        b"000000110000000001",b"000000111000000001",b"000001000000000001",b"000001001000000001",
        b"000001100000000001",b"000001101000000001",b"000001110000000001",b"000001111000000001",
        b"000010000000000001",b"000010001000000001",b"000010010000000001",b"000010011000000001",
        b"000010100000000001",b"000010101000000001",b"000010110000000001",b"000011000000000001",
        b"000011001000000001",b"000011010000000001",b"000011011000000001",b"000011100000000001",
        b"000011101000000001",b"000011110000000001",b"000011111000000001",b"000100000000000001",
        b"000100001000000001",b"000100010000000001",b"000100011000000001",b"000100100000000001",
        -- Row: 2
        b"000000001000000010",b"000000010000000010",b"000000011000000010",b"000000100000000010",
        b"000000111000000010",b"000001000000000010",b"000001001000000010",b"000001010000000010",
        b"000001011000000010",b"000001100000000010",b"000001101000000010",b"000001111000000010",
        b"000010000000000010",b"000010011000000010",b"000010100000000010",b"000010101000000010",
        b"000010110000000010",b"000010111000000010",b"000011000000000010",b"000011001000000010",
        b"000011011000000010",b"000011100000000010",b"000011101000000010",b"000011110000000010",
        b"000011111000000010",b"000100001000000010",b"000100010000000010",b"000100011000000010",
        b"000100100000000010",b"000100101000000010",b"000100110000000010",
        -- Row: 3
        b"000000001000000011",b"000000010000000011",b"000000011000000011",b"000000100000000011",
        b"000000101000000011",b"000000111000000011",b"000001000000000011",b"000001001000000011",
        b"000001010000000011",b"000001011000000011",b"000001100000000011",b"000001101000000011",
        b"000001110000000011",b"000001111000000011",b"000010000000000011",b"000010001000000011",
        b"000010011000000011",b"000010100000000011",b"000010110000000011",b"000010111000000011",
        b"000011000000000011",b"000011001000000011",b"000011010000000011",b"000011011000000011",
        b"000011101000000011",b"000011110000000011",b"000011111000000011",b"000100010000000011",
        b"000100011000000011",b"000100100000000011",b"000100101000000011",b"000100110000000011",
        -- Row: 4
        b"000000001000000100",b"000000010000000100",b"000000011000000100",b"000000100000000100",
        b"000000101000000100",b"000000110000000100",b"000000111000000100",b"000001000000000100",
        b"000001001000000100",b"000001010000000100",b"000001100000000100",b"000001101000000100",
        b"000001110000000100",b"000001111000000100",b"000010000000000100",b"000010010000000100",
        b"000010011000000100",b"000010100000000100",b"000010101000000100",b"000010110000000100",
        b"000010111000000100",b"000011000000000100",b"000011001000000100",b"000011010000000100",
        b"000011011000000100",b"000011100000000100",b"000011110000000100",b"000011111000000100",
        b"000100000000000100",b"000100001000000100",b"000100011000000100",b"000100100000000100",
        b"000100110000000100",
        -- Row: 5
        b"000000001000000101",b"000000011000000101",b"000000101000000101",b"000000110000000101",
        b"000000111000000101",b"000001001000000101",b"000001010000000101",b"000001011000000101",
        b"000001100000000101",b"000001101000000101",b"000001111000000101",b"000010000000000101",
        b"000010001000000101",b"000010010000000101",b"000010011000000101",b"000010100000000101",
        b"000010101000000101",b"000010110000000101",b"000010111000000101",b"000011000000000101",
        b"000011001000000101",b"000011010000000101",b"000011011000000101",b"000011101000000101",
        b"000011110000000101",b"000011111000000101",b"000100000000000101",b"000100001000000101",
        b"000100010000000101",b"000100011000000101",b"000100100000000101",b"000100110000000101",
        -- Row: 6
        b"000000001000000110",b"000000011000000110",b"000000100000000110",b"000000101000000110",
        b"000000110000000110",b"000000111000000110",b"000001000000000110",b"000001001000000110",
        b"000001011000000110",b"000001100000000110",b"000001111000000110",b"000010000000000110",
        b"000010001000000110",b"000010010000000110",b"000010011000000110",b"000010101000000110",
        b"000010110000000110",b"000010111000000110",b"000011011000000110",b"000011100000000110",
        b"000011101000000110",b"000011110000000110",b"000011111000000110",b"000100000000000110",
        b"000100001000000110",b"000100010000000110",b"000100011000000110",b"000100100000000110",
        b"000100101000000110",
        -- Row: 7
        b"000000001000000111",b"000000011000000111",b"000000100000000111",b"000000101000000111",
        b"000000111000000111",b"000001000000000111",b"000001001000000111",b"000001011000000111",
        b"000001100000000111",b"000001101000000111",b"000001110000000111",b"000001111000000111",
        b"000010000000000111",b"000010001000000111",b"000010010000000111",b"000010011000000111",
        b"000010100000000111",b"000010110000000111",b"000010111000000111",b"000011001000000111",
        b"000011010000000111",b"000011011000000111",b"000011100000000111",b"000011101000000111",
        b"000011110000000111",b"000011111000000111",b"000100010000000111",b"000100011000000111",
        b"000100100000000111",b"000100101000000111",b"000100110000000111",
        -- Row: 8
        b"000000001000001000",b"000000010000001000",b"000000011000001000",b"000000100000001000",
        b"000000111000001000",b"000001000000001000",b"000001001000001000",b"000001010000001000",
        b"000001011000001000",b"000001100000001000",b"000001101000001000",b"000001110000001000",
        b"000001111000001000",b"000010010000001000",b"000010011000001000",b"000010101000001000",
        b"000010110000001000",b"000010111000001000",b"000011001000001000",b"000011011000001000",
        b"000011100000001000",b"000011101000001000",b"000011110000001000",b"000011111000001000",
        b"000100000000001000",b"000100001000001000",b"000100010000001000",b"000100011000001000",
        b"000100100000001000",b"000100101000001000",b"000100110000001000",
        -- Row: 9
        b"000000001000001001",b"000000010000001001",b"000000011000001001",b"000000101000001001",
        b"000000110000001001",b"000000111000001001",b"000001000000001001",b"000001001000001001",
        b"000001010000001001",b"000001011000001001",b"000001101000001001",b"000001110000001001",
        b"000001111000001001",b"000010001000001001",b"000010010000001001",b"000010011000001001",
        b"000010100000001001",b"000010101000001001",b"000010110000001001",b"000010111000001001",
        b"000011000000001001",b"000011001000001001",b"000011010000001001",b"000011011000001001",
        b"000011100000001001",b"000011101000001001",b"000011110000001001",b"000011111000001001",
        b"000100000000001001",b"000100001000001001",b"000100011000001001",b"000100100000001001",
        b"000100101000001001",b"000100110000001001",
        -- Row: 10
        b"000000001000001010",b"000000010000001010",b"000000011000001010",b"000000100000001010",
        b"000000101000001010",b"000000110000001010",b"000000111000001010",b"000001000000001010",
        b"000001010000001010",b"000001011000001010",b"000001101000001010",b"000001110000001010",
        b"000001111000001010",b"000010000000001010",b"000010001000001010",b"000010010000001010",
        b"000010100000001010",b"000010101000001010",b"000010111000001010",b"000011000000001010",
        b"000011001000001010",b"000011010000001010",b"000011011000001010",b"000011100000001010",
        b"000011110000001010",b"000011111000001010",b"000100000000001010",b"000100011000001010",
        b"000100100000001010",b"000100101000001010",b"000100110000001010",
        -- Row: 11
        b"000000001000001011",b"000000011000001011",b"000000100000001011",b"000000101000001011",
        b"000000110000001011",b"000000111000001011",b"000001000000001011",b"000001001000001011",
        b"000001010000001011",b"000001011000001011",b"000001100000001011",b"000001110000001011",
        b"000001111000001011",b"000010000000001011",b"000010001000001011",b"000010010000001011",
        b"000010011000001011",b"000010101000001011",b"000010110000001011",b"000011000000001011",
        b"000011001000001011",b"000011010000001011",b"000011011000001011",b"000011100000001011",
        b"000011110000001011",b"000100000000001011",b"000100001000001011",b"000100010000001011",
        b"000100011000001011",b"000100100000001011",b"000100101000001011",b"000100110000001011",
        -- Row: 12
        b"000000001000001100",b"000000010000001100",b"000000011000001100",b"000000100000001100",
        b"000000101000001100",b"000000110000001100",b"000000111000001100",b"000001000000001100",
        b"000001001000001100",b"000001010000001100",b"000001011000001100",b"000001100000001100",
        b"000001101000001100",b"000001110000001100",b"000001111000001100",b"000010000000001100",
        b"000010001000001100",b"000010010000001100",b"000010011000001100",b"000010100000001100",
        b"000010101000001100",b"000010110000001100",b"000010111000001100",b"000011000000001100",
        b"000011001000001100",b"000011010000001100",b"000011011000001100",b"000011100000001100",
        b"000011101000001100",b"000011111000001100",b"000100000000001100",b"000100001000001100",
        b"000100010000001100",b"000100011000001100",b"000100100000001100",b"000100101000001100",
        -- Row: 13
        b"000000001000001101",b"000000010000001101",b"000000011000001101",b"000000100000001101",
        b"000000101000001101",b"000000110000001101",b"000000111000001101",b"000001000000001101",
        b"000001001000001101",b"000001010000001101",b"000001011000001101",b"000001100000001101",
        b"000001110000001101",b"000001111000001101",b"000010000000001101",b"000010001000001101",
        b"000010011000001101",b"000010100000001101",b"000010101000001101",b"000010110000001101",
        b"000010111000001101",b"000011000000001101",b"000011001000001101",b"000011011000001101",
        b"000011100000001101",b"000011101000001101",b"000011110000001101",b"000011111000001101",
        b"000100000000001101",b"000100001000001101",b"000100010000001101",b"000100011000001101",
        b"000100100000001101",b"000100101000001101",
        -- Row: 14
        b"000000001000001110",b"000000101000001110",b"000000110000001110",b"000000111000001110",
        b"000001010000001110",b"000001011000001110",b"000001100000001110",b"000001101000001110",
        b"000001110000001110",b"000001111000001110",b"000010000000001110",b"000010001000001110",
        b"000010010000001110",b"000010011000001110",b"000010100000001110",b"000010101000001110",
        b"000010110000001110",b"000010111000001110",b"000011000000001110",b"000011001000001110",
        b"000011011000001110",b"000011100000001110",b"000011101000001110",b"000011110000001110",
        b"000011111000001110",b"000100000000001110",b"000100011000001110",b"000100100000001110",
        b"000100101000001110",b"000100110000001110",
        -- Row: 15
        b"000000001000001111",b"000000010000001111",b"000000011000001111",b"000000101000001111",
        b"000000110000001111",b"000001001000001111",b"000001010000001111",b"000001100000001111",
        b"000001101000001111",b"000001110000001111",b"000001111000001111",b"000010010000001111",
        b"000010011000001111",b"000010100000001111",b"000010110000001111",b"000010111000001111",
        b"000011000000001111",b"000011010000001111",b"000011011000001111",b"000011100000001111",
        b"000011101000001111",b"000011110000001111",b"000011111000001111",b"000100000000001111",
        b"000100010000001111",b"000100011000001111",b"000100100000001111",b"000100101000001111",
        b"000100110000001111",
        -- Row: 16
        b"000000001000010000",b"000000010000010000",b"000000011000010000",b"000000101000010000",
        b"000000110000010000",b"000000111000010000",b"000001001000010000",b"000001010000010000",
        b"000001100000010000",b"000001101000010000",b"000001110000010000",b"000001111000010000",
        b"000010001000010000",b"000010010000010000",b"000010011000010000",b"000010100000010000",
        b"000010111000010000",b"000011001000010000",b"000011010000010000",b"000011011000010000",
        b"000011110000010000",b"000011111000010000",b"000100000000010000",b"000100001000010000",
        b"000100010000010000",b"000100011000010000",b"000100100000010000",b"000100101000010000",
        b"000100110000010000",
        -- Row: 17
        b"000000001000010001",b"000000010000010001",b"000000011000010001",b"000000100000010001",
        b"000000101000010001",b"000000110000010001",b"000000111000010001",b"000001001000010001",
        b"000001010000010001",b"000001011000010001",b"000001101000010001",b"000001111000010001",
        b"000010000000010001",b"000010001000010001",b"000010010000010001",b"000010011000010001",
        b"000010100000010001",b"000010110000010001",b"000010111000010001",b"000011000000010001",
        b"000011001000010001",b"000011010000010001",b"000011011000010001",b"000011101000010001",
        b"000011110000010001",b"000100000000010001",b"000100001000010001",b"000100010000010001",
        b"000100011000010001",b"000100100000010001",b"000100101000010001",
        -- Row: 18
        b"000000001000010010",b"000000010000010010",b"000000011000010010",b"000000100000010010",
        b"000000101000010010",b"000000110000010010",b"000000111000010010",b"000001000000010010",
        b"000001001000010010",b"000001010000010010",b"000001011000010010",b"000001100000010010",
        b"000001101000010010",b"000001110000010010",b"000001111000010010",b"000010000000010010",
        b"000010001000010010",b"000010010000010010",b"000010011000010010",b"000010110000010010",
        b"000010111000010010",b"000011000000010010",b"000011001000010010",b"000011010000010010",
        b"000011100000010010",b"000011101000010010",b"000011110000010010",b"000011111000010010",
        b"000100010000010010",b"000100011000010010",b"000100100000010010",b"000100101000010010",
        b"000100110000010010",
        -- Row: 19
        b"000000001000010011",b"000000010000010011",b"000000100000010011",b"000000101000010011",
        b"000000110000010011",b"000000111000010011",b"000001000000010011",b"000001001000010011",
        b"000001010000010011",b"000001011000010011",b"000001100000010011",b"000001101000010011",
        b"000001110000010011",b"000001111000010011",b"000010000000010011",b"000010010000010011",
        b"000010011000010011",b"000010100000010011",b"000010110000010011",b"000010111000010011",
        b"000011000000010011",b"000011001000010011",b"000011010000010011",b"000011011000010011",
        b"000011100000010011",b"000011101000010011",b"000011110000010011",b"000011111000010011",
        b"000100000000010011",b"000100010000010011",b"000100011000010011",b"000100100000010011",
        b"000100101000010011",b"000100110000010011",
        -- Row: 20
        b"000000001000010100",b"000000010000010100",b"000000011000010100",b"000000100000010100",
        b"000000101000010100",b"000000110000010100",b"000000111000010100",b"000001000000010100",
        b"000001001000010100",b"000001010000010100",b"000001011000010100",b"000001100000010100",
        b"000001101000010100",b"000001111000010100",b"000010000000010100",b"000010001000010100",
        b"000010010000010100",b"000010011000010100",b"000010100000010100",b"000010101000010100",
        b"000010111000010100",b"000011000000010100",b"000011001000010100",b"000011010000010100",
        b"000011011000010100",b"000011100000010100",b"000011101000010100",b"000011111000010100",
        b"000100000000010100",b"000100010000010100",b"000100011000010100",b"000100100000010100",
        b"000100101000010100",b"000100110000010100",
        -- Row: 21
        b"000000001000010101",b"000000010000010101",b"000000011000010101",b"000000100000010101",
        b"000000101000010101",b"000000111000010101",b"000001000000010101",b"000001001000010101",
        b"000001011000010101",b"000001100000010101",b"000001111000010101",b"000010000000010101",
        b"000010001000010101",b"000010010000010101",b"000010011000010101",b"000010100000010101",
        b"000010101000010101",b"000010110000010101",b"000010111000010101",b"000011000000010101",
        b"000011010000010101",b"000011011000010101",b"000011100000010101",b"000011101000010101",
        b"000011110000010101",b"000011111000010101",b"000100000000010101",b"000100001000010101",
        b"000100010000010101",b"000100011000010101",b"000100100000010101",b"000100101000010101",
        b"000100110000010101",
        -- Row: 22
        b"000000010000010110",b"000000011000010110",b"000000100000010110",b"000000101000010110",
        b"000000110000010110",b"000001000000010110",b"000001001000010110",b"000001010000010110",
        b"000001011000010110",b"000001100000010110",b"000001110000010110",b"000001111000010110",
        b"000010000000010110",b"000010001000010110",b"000010010000010110",b"000010100000010110",
        b"000010101000010110",b"000010110000010110",b"000010111000010110",b"000011001000010110",
        b"000011010000010110",b"000011011000010110",b"000011101000010110",b"000011110000010110",
        b"000011111000010110",b"000100000000010110",b"000100001000010110",b"000100010000010110",
        b"000100011000010110",b"000100100000010110",b"000100101000010110",
        -- Row: 23
        b"000000010000010111",b"000000011000010111",b"000000100000010111",b"000000110000010111",
        b"000000111000010111",b"000001000000010111",b"000001001000010111",b"000001010000010111",
        b"000001011000010111",b"000001100000010111",b"000001110000010111",b"000001111000010111",
        b"000010000000010111",b"000010011000010111",b"000010100000010111",b"000010101000010111",
        b"000010110000010111",b"000010111000010111",b"000011001000010111",b"000011010000010111",
        b"000011011000010111",b"000011110000010111",b"000011111000010111",b"000100000000010111",
        b"000100001000010111",b"000100011000010111",b"000100100000010111",b"000100101000010111",
        b"000100110000010111",
        -- Row: 24
        b"000000001000011000",b"000000010000011000",b"000000101000011000",b"000000110000011000",
        b"000000111000011000",b"000001000000011000",b"000001001000011000",b"000001010000011000",
        b"000001011000011000",b"000001100000011000",b"000001101000011000",b"000001110000011000",
        b"000001111000011000",b"000010000000011000",b"000010001000011000",b"000010010000011000",
        b"000010011000011000",b"000010100000011000",b"000010101000011000",b"000010110000011000",
        b"000010111000011000",b"000011000000011000",b"000011001000011000",b"000011010000011000",
        b"000011011000011000",b"000011100000011000",b"000011101000011000",b"000011111000011000",
        b"000100000000011000",b"000100010000011000",b"000100100000011000",b"000100101000011000",
        b"000100110000011000",
        -- Row: 25
        b"000000001000011001",b"000000010000011001",b"000000011000011001",b"000000101000011001",
        b"000000110000011001",b"000000111000011001",b"000001000000011001",b"000001001000011001",
        b"000001010000011001",b"000001100000011001",b"000001101000011001",b"000001110000011001",
        b"000001111000011001",b"000010000000011001",b"000010001000011001",b"000010010000011001",
        b"000010011000011001",b"000010100000011001",b"000010101000011001",b"000010110000011001",
        b"000010111000011001",b"000011000000011001",b"000011010000011001",b"000011011000011001",
        b"000011110000011001",b"000011111000011001",b"000100000000011001",b"000100001000011001",
        b"000100010000011001",b"000100011000011001",b"000100100000011001",b"000100101000011001",
        b"000100110000011001",
        -- Row: 26
        b"000000001000011010",b"000000010000011010",b"000000011000011010",b"000000100000011010",
        b"000000101000011010",b"000000110000011010",b"000001000000011010",b"000001001000011010",
        b"000001011000011010",b"000001100000011010",b"000001101000011010",b"000001110000011010",
        b"000010000000011010",b"000010001000011010",b"000010010000011010",b"000010100000011010",
        b"000010110000011010",b"000010111000011010",b"000011000000011010",b"000011001000011010",
        b"000011010000011010",b"000011011000011010",b"000011100000011010",b"000011101000011010",
        b"000011110000011010",b"000011111000011010",b"000100000000011010",b"000100001000011010",
        b"000100010000011010",b"000100011000011010",b"000100100000011010",b"000100110000011010",
        -- Row: 27
        b"000000001000011011",b"000000011000011011",b"000000100000011011",b"000000101000011011",
        b"000000111000011011",b"000001000000011011",b"000001001000011011",b"000001010000011011",
        b"000001011000011011",b"000001100000011011",b"000001101000011011",b"000001111000011011",
        b"000010000000011011",b"000010001000011011",b"000010100000011011",b"000010101000011011",
        b"000010110000011011",b"000010111000011011",b"000011000000011011",b"000011001000011011",
        b"000011010000011011",b"000011011000011011",b"000011100000011011",b"000011101000011011",
        b"000011110000011011",b"000100001000011011",b"000100010000011011",b"000100011000011011",
        b"000100110000011011",
        -- Row: 28
        b"000000010000011100",b"000000011000011100",b"000000100000011100",b"000001000000011100",
        b"000001001000011100",b"000001010000011100",b"000001011000011100",b"000001100000011100",
        b"000001101000011100",b"000001110000011100",b"000001111000011100",b"000010000000011100",
        b"000010011000011100",b"000010100000011100",b"000010101000011100",b"000010110000011100",
        b"000010111000011100",b"000011000000011100",b"000011001000011100",b"000011010000011100",
        b"000011011000011100",b"000011100000011100",b"000011101000011100",b"000100000000011100",
        b"000100001000011100",b"000100010000011100",b"000100011000011100",b"000100100000011100",
        b"000100101000011100"
        -- Row: 29
	    );
	
	type track_3_free_pos_mem_t is array (0 to 932) of signed(17 downto 0);
	constant track_3_free_pos_mem_c : track_3_free_pos_mem_t := (
        -- Row: 0
        -- Row: 1
        b"000000010000000001",b"000000100000000001",b"000000101000000001",b"000000110000000001",
        b"000000111000000001",b"000001000000000001",b"000001001000000001",b"000001011000000001",
        b"000001100000000001",b"000001101000000001",b"000001110000000001",b"000001111000000001",
        b"000010000000000001",b"000010001000000001",b"000010010000000001",b"000010011000000001",
        b"000010100000000001",b"000010110000000001",b"000010111000000001",b"000011000000000001",
        b"000011001000000001",b"000011010000000001",b"000011100000000001",b"000011101000000001",
        b"000011110000000001",b"000011111000000001",b"000100001000000001",b"000100010000000001",
        b"000100011000000001",
        -- Row: 2
        b"000000001000000010",b"000000010000000010",b"000000011000000010",b"000000100000000010",
        b"000000101000000010",b"000000110000000010",b"000000111000000010",b"000001000000000010",
        b"000001001000000010",b"000001010000000010",b"000001011000000010",b"000001100000000010",
        b"000001101000000010",b"000001110000000010",b"000001111000000010",b"000010001000000010",
        b"000010010000000010",b"000010011000000010",b"000010100000000010",b"000010101000000010",
        b"000010110000000010",b"000011000000000010",b"000011001000000010",b"000011010000000010",
        b"000011011000000010",b"000011100000000010",b"000011101000000010",b"000011110000000010",
        b"000011111000000010",b"000100000000000010",b"000100001000000010",b"000100010000000010",
        b"000100011000000010",b"000100100000000010",b"000100110000000010",
        -- Row: 3
        b"000000001000000011",b"000000010000000011",b"000000011000000011",b"000000100000000011",
        b"000000101000000011",b"000000110000000011",b"000001000000000011",b"000001001000000011",
        b"000001010000000011",b"000001011000000011",b"000001100000000011",b"000001101000000011",
        b"000001110000000011",b"000001111000000011",b"000010000000000011",b"000010010000000011",
        b"000010100000000011",b"000010101000000011",b"000010110000000011",b"000010111000000011",
        b"000011000000000011",b"000011001000000011",b"000011010000000011",b"000011011000000011",
        b"000011100000000011",b"000011101000000011",b"000011110000000011",b"000011111000000011",
        b"000100000000000011",b"000100001000000011",b"000100010000000011",b"000100011000000011",
        b"000100100000000011",b"000100101000000011",b"000100110000000011",
        -- Row: 4
        b"000000001000000100",b"000000010000000100",b"000000011000000100",b"000000100000000100",
        b"000000101000000100",b"000000110000000100",b"000000111000000100",b"000001000000000100",
        b"000001001000000100",b"000001010000000100",b"000001011000000100",b"000001100000000100",
        b"000001101000000100",b"000001110000000100",b"000001111000000100",b"000010000000000100",
        b"000010001000000100",b"000010011000000100",b"000010100000000100",b"000010101000000100",
        b"000010110000000100",b"000010111000000100",b"000011000000000100",b"000011001000000100",
        b"000011010000000100",b"000011011000000100",b"000011100000000100",b"000011101000000100",
        b"000011111000000100",b"000100000000000100",b"000100001000000100",b"000100010000000100",
        b"000100011000000100",b"000100100000000100",b"000100101000000100",b"000100110000000100",
        -- Row: 5
        b"000000001000000101",b"000000010000000101",b"000000100000000101",b"000000101000000101",
        b"000000110000000101",b"000000111000000101",b"000001000000000101",b"000001001000000101",
        b"000001010000000101",b"000001100000000101",b"000001101000000101",b"000001110000000101",
        b"000001111000000101",b"000010000000000101",b"000010001000000101",b"000010010000000101",
        b"000010011000000101",b"000010100000000101",b"000010101000000101",b"000010110000000101",
        b"000010111000000101",b"000011000000000101",b"000011001000000101",b"000011010000000101",
        b"000011011000000101",b"000011101000000101",b"000011110000000101",b"000011111000000101",
        b"000100000000000101",b"000100010000000101",b"000100011000000101",b"000100100000000101",
        b"000100101000000101",b"000100110000000101",
        -- Row: 6
        b"000000001000000110",b"000000010000000110",b"000000011000000110",b"000000100000000110",
        b"000000101000000110",b"000000110000000110",b"000000111000000110",b"000001000000000110",
        b"000001001000000110",b"000001010000000110",b"000001011000000110",b"000001100000000110",
        b"000001101000000110",b"000001110000000110",b"000001111000000110",b"000010000000000110",
        b"000010001000000110",b"000010010000000110",b"000010011000000110",b"000010100000000110",
        b"000010101000000110",b"000010110000000110",b"000011000000000110",b"000011001000000110",
        b"000011010000000110",b"000011100000000110",b"000011101000000110",b"000011110000000110",
        b"000011111000000110",b"000100000000000110",b"000100011000000110",b"000100100000000110",
        b"000100101000000110",b"000100110000000110",
        -- Row: 7
        b"000000010000000111",b"000000011000000111",b"000000100000000111",b"000000110000000111",
        b"000000111000000111",b"000001001000000111",b"000001010000000111",b"000001011000000111",
        b"000001100000000111",b"000001101000000111",b"000001110000000111",b"000001111000000111",
        b"000010000000000111",b"000010001000000111",b"000010010000000111",b"000010011000000111",
        b"000010100000000111",b"000010101000000111",b"000010110000000111",b"000010111000000111",
        b"000011000000000111",b"000011001000000111",b"000011010000000111",b"000011011000000111",
        b"000011100000000111",b"000011101000000111",b"000011110000000111",b"000011111000000111",
        b"000100001000000111",b"000100010000000111",b"000100011000000111",b"000100100000000111",
        b"000100101000000111",
        -- Row: 8
        b"000000010000001000",b"000000011000001000",b"000000100000001000",b"000000110000001000",
        b"000001000000001000",b"000001001000001000",b"000001010000001000",b"000001011000001000",
        b"000001100000001000",b"000001110000001000",b"000001111000001000",b"000010000000001000",
        b"000010010000001000",b"000010011000001000",b"000010100000001000",b"000010101000001000",
        b"000010110000001000",b"000010111000001000",b"000011000000001000",b"000011001000001000",
        b"000011010000001000",b"000011011000001000",b"000011100000001000",b"000011101000001000",
        b"000011110000001000",b"000011111000001000",b"000100000000001000",b"000100001000001000",
        b"000100010000001000",b"000100011000001000",b"000100100000001000",b"000100101000001000",
        -- Row: 9
        b"000000001000001001",b"000000010000001001",b"000000011000001001",b"000000100000001001",
        b"000000101000001001",b"000000110000001001",b"000001000000001001",b"000001001000001001",
        b"000001010000001001",b"000001011000001001",b"000001101000001001",b"000001110000001001",
        b"000001111000001001",b"000010001000001001",b"000010010000001001",b"000010011000001001",
        b"000010101000001001",b"000010110000001001",b"000011000000001001",b"000011001000001001",
        b"000011010000001001",b"000011011000001001",b"000011100000001001",b"000011101000001001",
        b"000011110000001001",b"000011111000001001",b"000100000000001001",b"000100001000001001",
        b"000100011000001001",b"000100100000001001",b"000100101000001001",b"000100110000001001",
        -- Row: 10
        b"000000001000001010",b"000000010000001010",b"000000011000001010",b"000000100000001010",
        b"000000101000001010",b"000000110000001010",b"000000111000001010",b"000001000000001010",
        b"000001001000001010",b"000001010000001010",b"000001011000001010",b"000001100000001010",
        b"000001110000001010",b"000001111000001010",b"000010001000001010",b"000010010000001010",
        b"000010011000001010",b"000010111000001010",b"000011000000001010",b"000011001000001010",
        b"000011010000001010",b"000011011000001010",b"000011100000001010",b"000011101000001010",
        b"000011110000001010",b"000011111000001010",b"000100000000001010",b"000100001000001010",
        b"000100010000001010",b"000100011000001010",b"000100100000001010",b"000100101000001010",
        b"000100110000001010",
        -- Row: 11
        b"000000001000001011",b"000000010000001011",b"000000100000001011",b"000000101000001011",
        b"000000110000001011",b"000000111000001011",b"000001000000001011",b"000001001000001011",
        b"000001010000001011",b"000001011000001011",b"000001100000001011",b"000001101000001011",
        b"000001110000001011",b"000001111000001011",b"000010000000001011",b"000010001000001011",
        b"000010010000001011",b"000010011000001011",b"000010100000001011",b"000010101000001011",
        b"000010110000001011",b"000010111000001011",b"000011000000001011",b"000011001000001011",
        b"000011010000001011",b"000011011000001011",b"000011100000001011",b"000011110000001011",
        b"000011111000001011",b"000100000000001011",b"000100001000001011",b"000100010000001011",
        b"000100011000001011",b"000100100000001011",b"000100101000001011",b"000100110000001011",
        -- Row: 12
        b"000000001000001100",b"000000010000001100",b"000000011000001100",b"000000100000001100",
        b"000000101000001100",b"000000110000001100",b"000000111000001100",b"000001000000001100",
        b"000001010000001100",b"000001011000001100",b"000001100000001100",b"000001101000001100",
        b"000001110000001100",b"000001111000001100",b"000010000000001100",b"000010001000001100",
        b"000010010000001100",b"000010011000001100",b"000010100000001100",b"000010101000001100",
        b"000010110000001100",b"000010111000001100",b"000011000000001100",b"000011001000001100",
        b"000011010000001100",b"000011101000001100",b"000011110000001100",b"000011111000001100",
        b"000100000000001100",b"000100001000001100",b"000100010000001100",b"000100011000001100",
        b"000100101000001100",b"000100110000001100",
        -- Row: 13
        b"000000010000001101",b"000000011000001101",b"000000100000001101",b"000000101000001101",
        b"000000110000001101",b"000000111000001101",b"000001000000001101",b"000001011000001101",
        b"000001100000001101",b"000001101000001101",b"000001110000001101",b"000001111000001101",
        b"000010000000001101",b"000010001000001101",b"000010010000001101",b"000010011000001101",
        b"000010100000001101",b"000010101000001101",b"000010110000001101",b"000010111000001101",
        b"000011000000001101",b"000011001000001101",b"000011010000001101",b"000011011000001101",
        b"000011100000001101",b"000011101000001101",b"000011110000001101",b"000011111000001101",
        b"000100001000001101",b"000100010000001101",b"000100011000001101",b"000100100000001101",
        b"000100110000001101",
        -- Row: 14
        b"000000010000001110",b"000000011000001110",b"000000100000001110",b"000000101000001110",
        b"000000111000001110",b"000001000000001110",b"000001001000001110",b"000001010000001110",
        b"000001011000001110",b"000001100000001110",b"000001101000001110",b"000001110000001110",
        b"000010000000001110",b"000010001000001110",b"000010011000001110",b"000010100000001110",
        b"000010101000001110",b"000010110000001110",b"000010111000001110",b"000011000000001110",
        b"000011001000001110",b"000011010000001110",b"000011011000001110",b"000011100000001110",
        b"000011101000001110",b"000011110000001110",b"000100000000001110",b"000100001000001110",
        b"000100010000001110",b"000100011000001110",b"000100100000001110",b"000100110000001110",
        -- Row: 15
        b"000000001000001111",b"000000011000001111",b"000000100000001111",b"000000101000001111",
        b"000000110000001111",b"000001000000001111",b"000001001000001111",b"000001010000001111",
        b"000001011000001111",b"000001100000001111",b"000001101000001111",b"000001110000001111",
        b"000001111000001111",b"000010000000001111",b"000010010000001111",b"000010100000001111",
        b"000010101000001111",b"000010110000001111",b"000011000000001111",b"000011001000001111",
        b"000011010000001111",b"000011011000001111",b"000011100000001111",b"000011101000001111",
        b"000011110000001111",b"000011111000001111",b"000100001000001111",b"000100010000001111",
        b"000100011000001111",b"000100100000001111",b"000100101000001111",
        -- Row: 16
        b"000000001000010000",b"000000010000010000",b"000000011000010000",b"000000100000010000",
        b"000000101000010000",b"000000110000010000",b"000001000000010000",b"000001001000010000",
        b"000001010000010000",b"000001011000010000",b"000001100000010000",b"000001101000010000",
        b"000001110000010000",b"000001111000010000",b"000010000000010000",b"000010001000010000",
        b"000010010000010000",b"000010011000010000",b"000010100000010000",b"000010101000010000",
        b"000010111000010000",b"000011001000010000",b"000011010000010000",b"000011011000010000",
        b"000011100000010000",b"000011101000010000",b"000011110000010000",b"000011111000010000",
        b"000100000000010000",b"000100001000010000",b"000100010000010000",b"000100011000010000",
        b"000100100000010000",b"000100101000010000",b"000100110000010000",
        -- Row: 17
        b"000000001000010001",b"000000010000010001",b"000000011000010001",b"000000100000010001",
        b"000000101000010001",b"000000110000010001",b"000000111000010001",b"000001000000010001",
        b"000001001000010001",b"000001010000010001",b"000001011000010001",b"000001100000010001",
        b"000001101000010001",b"000001110000010001",b"000001111000010001",b"000010000000010001",
        b"000010001000010001",b"000010010000010001",b"000010011000010001",b"000010100000010001",
        b"000010101000010001",b"000010110000010001",b"000010111000010001",b"000011000000010001",
        b"000011001000010001",b"000011011000010001",b"000011100000010001",b"000011101000010001",
        b"000011110000010001",b"000011111000010001",b"000100000000010001",b"000100001000010001",
        b"000100010000010001",b"000100011000010001",b"000100100000010001",b"000100101000010001",
        b"000100110000010001",
        -- Row: 18
        b"000000001000010010",b"000000011000010010",b"000000100000010010",b"000000101000010010",
        b"000000110000010010",b"000000111000010010",b"000001000000010010",b"000001001000010010",
        b"000001010000010010",b"000001011000010010",b"000001100000010010",b"000001111000010010",
        b"000010000000010010",b"000010001000010010",b"000010010000010010",b"000010011000010010",
        b"000010100000010010",b"000010101000010010",b"000010110000010010",b"000010111000010010",
        b"000011000000010010",b"000011001000010010",b"000011010000010010",b"000011011000010010",
        b"000011100000010010",b"000011101000010010",b"000011110000010010",b"000011111000010010",
        b"000100000000010010",b"000100001000010010",b"000100010000010010",b"000100011000010010",
        b"000100100000010010",b"000100101000010010",b"000100110000010010",
        -- Row: 19
        b"000000001000010011",b"000000011000010011",b"000000100000010011",b"000000110000010011",
        b"000000111000010011",b"000001000000010011",b"000001001000010011",b"000001010000010011",
        b"000001011000010011",b"000001100000010011",b"000001101000010011",b"000001111000010011",
        b"000010000000010011",b"000010001000010011",b"000010011000010011",b"000010100000010011",
        b"000010101000010011",b"000010110000010011",b"000010111000010011",b"000011000000010011",
        b"000011001000010011",b"000011010000010011",b"000011011000010011",b"000011100000010011",
        b"000011110000010011",b"000011111000010011",b"000100000000010011",b"000100001000010011",
        b"000100010000010011",b"000100011000010011",b"000100100000010011",b"000100101000010011",
        b"000100110000010011",
        -- Row: 20
        b"000000001000010100",b"000000010000010100",b"000000100000010100",b"000000101000010100",
        b"000000110000010100",b"000000111000010100",b"000001000000010100",b"000001011000010100",
        b"000001100000010100",b"000001101000010100",b"000001111000010100",b"000010000000010100",
        b"000010001000010100",b"000010010000010100",b"000010011000010100",b"000010101000010100",
        b"000010110000010100",b"000010111000010100",b"000011000000010100",b"000011001000010100",
        b"000011010000010100",b"000011011000010100",b"000011110000010100",b"000011111000010100",
        b"000100000000010100",b"000100011000010100",b"000100110000010100",
        -- Row: 21
        b"000000001000010101",b"000000010000010101",b"000000011000010101",b"000000100000010101",
        b"000000101000010101",b"000000110000010101",b"000000111000010101",b"000001000000010101",
        b"000001001000010101",b"000001011000010101",b"000001100000010101",b"000001101000010101",
        b"000001110000010101",b"000001111000010101",b"000010000000010101",b"000010001000010101",
        b"000010010000010101",b"000010011000010101",b"000010100000010101",b"000010101000010101",
        b"000010110000010101",b"000010111000010101",b"000011000000010101",b"000011001000010101",
        b"000011010000010101",b"000011011000010101",b"000011100000010101",b"000011101000010101",
        b"000011110000010101",b"000011111000010101",b"000100000000010101",b"000100010000010101",
        b"000100011000010101",b"000100101000010101",b"000100110000010101",
        -- Row: 22
        b"000000001000010110",b"000000010000010110",b"000000011000010110",b"000000100000010110",
        b"000000101000010110",b"000000110000010110",b"000000111000010110",b"000001000000010110",
        b"000001001000010110",b"000001010000010110",b"000001011000010110",b"000001100000010110",
        b"000001101000010110",b"000001110000010110",b"000001111000010110",b"000010000000010110",
        b"000010001000010110",b"000010010000010110",b"000010011000010110",b"000010100000010110",
        b"000010101000010110",b"000010110000010110",b"000010111000010110",b"000011001000010110",
        b"000011010000010110",b"000011011000010110",b"000011100000010110",b"000011101000010110",
        b"000011110000010110",b"000011111000010110",b"000100001000010110",b"000100010000010110",
        b"000100011000010110",b"000100100000010110",b"000100110000010110",
        -- Row: 23
        b"000000001000010111",b"000000010000010111",b"000000011000010111",b"000000101000010111",
        b"000000110000010111",b"000000111000010111",b"000001000000010111",b"000001001000010111",
        b"000001010000010111",b"000001011000010111",b"000001100000010111",b"000001110000010111",
        b"000001111000010111",b"000010000000010111",b"000010001000010111",b"000010010000010111",
        b"000010011000010111",b"000010100000010111",b"000010101000010111",b"000010110000010111",
        b"000010111000010111",b"000011010000010111",b"000011011000010111",b"000011100000010111",
        b"000011101000010111",b"000011110000010111",b"000011111000010111",b"000100000000010111",
        b"000100001000010111",b"000100010000010111",b"000100011000010111",b"000100100000010111",
        b"000100101000010111",b"000100110000010111",
        -- Row: 24
        b"000000001000011000",b"000000010000011000",b"000000011000011000",b"000000101000011000",
        b"000000110000011000",b"000000111000011000",b"000001000000011000",b"000001001000011000",
        b"000001010000011000",b"000001011000011000",b"000001101000011000",b"000001110000011000",
        b"000001111000011000",b"000010000000011000",b"000010010000011000",b"000010100000011000",
        b"000010101000011000",b"000010110000011000",b"000010111000011000",b"000011000000011000",
        b"000011001000011000",b"000011010000011000",b"000011011000011000",b"000011100000011000",
        b"000011110000011000",b"000011111000011000",b"000100000000011000",b"000100001000011000",
        b"000100010000011000",b"000100011000011000",b"000100100000011000",b"000100101000011000",
        b"000100110000011000",
        -- Row: 25
        b"000000001000011001",b"000000010000011001",b"000000011000011001",b"000000100000011001",
        b"000000101000011001",b"000000110000011001",b"000001000000011001",b"000001001000011001",
        b"000001010000011001",b"000001011000011001",b"000001100000011001",b"000001101000011001",
        b"000001110000011001",b"000001111000011001",b"000010000000011001",b"000010001000011001",
        b"000010100000011001",b"000010101000011001",b"000010110000011001",b"000010111000011001",
        b"000011000000011001",b"000011001000011001",b"000011010000011001",b"000011011000011001",
        b"000011100000011001",b"000011101000011001",b"000011110000011001",b"000011111000011001",
        b"000100000000011001",b"000100010000011001",b"000100011000011001",b"000100100000011001",
        b"000100101000011001",b"000100110000011001",
        -- Row: 26
        b"000000010000011010",b"000000011000011010",b"000000100000011010",b"000000101000011010",
        b"000000110000011010",b"000000111000011010",b"000001000000011010",b"000001001000011010",
        b"000001010000011010",b"000001011000011010",b"000001100000011010",b"000001101000011010",
        b"000001110000011010",b"000010000000011010",b"000010001000011010",b"000010010000011010",
        b"000010011000011010",b"000010100000011010",b"000010101000011010",b"000010110000011010",
        b"000011000000011010",b"000011001000011010",b"000011010000011010",b"000011011000011010",
        b"000011100000011010",b"000011101000011010",b"000011110000011010",b"000011111000011010",
        b"000100000000011010",b"000100001000011010",b"000100010000011010",b"000100011000011010",
        b"000100101000011010",b"000100110000011010",
        -- Row: 27
        b"000000010000011011",b"000000011000011011",b"000000100000011011",b"000000101000011011",
        b"000000110000011011",b"000000111000011011",b"000001001000011011",b"000001010000011011",
        b"000001011000011011",b"000001100000011011",b"000001101000011011",b"000001111000011011",
        b"000010000000011011",b"000010001000011011",b"000010010000011011",b"000010011000011011",
        b"000010100000011011",b"000010101000011011",b"000010111000011011",b"000011000000011011",
        b"000011001000011011",b"000011010000011011",b"000011011000011011",b"000011100000011011",
        b"000011101000011011",b"000011110000011011",b"000011111000011011",b"000100000000011011",
        b"000100001000011011",b"000100010000011011",b"000100011000011011",b"000100100000011011",
        b"000100110000011011",
        -- Row: 28
        b"000000011000011100",b"000000100000011100",b"000000101000011100",b"000000110000011100",
        b"000001010000011100",b"000001011000011100",b"000001100000011100",b"000001101000011100",
        b"000001111000011100",b"000010000000011100",b"000010001000011100",b"000010010000011100",
        b"000010011000011100",b"000010100000011100",b"000010101000011100",b"000010110000011100",
        b"000010111000011100",b"000011000000011100",b"000011001000011100",b"000011010000011100",
        b"000011011000011100",b"000011100000011100",b"000011111000011100",b"000100000000011100",
        b"000100001000011100",b"000100011000011100",b"000100100000011100",b"000100101000011100",
        b"000100110000011100"
        -- Row: 29
	);
	
	type track_4_free_pos_mem_t is array (0 to 660) of signed(17 downto 0);
	constant track_4_free_pos_mem_c : track_4_free_pos_mem_t := (
	
        -- Row: 0
        -- Row: 1
        b"000000010000000001",b"000000011000000001",b"000000100000000001",b"000000101000000001",
        b"000000110000000001",b"000000111000000001",b"000001000000000001",b"000001001000000001",
        b"000001010000000001",b"000001011000000001",b"000001111000000001",b"000010000000000001",
        b"000010001000000001",b"000010010000000001",b"000010011000000001",b"000010110000000001",
        b"000010111000000001",b"000011000000000001",b"000011001000000001",b"000011010000000001",
        b"000011011000000001",b"000011100000000001",b"000011101000000001",b"000011110000000001",
        b"000011111000000001",b"000100000000000001",b"000100001000000001",b"000100010000000001",
        b"000100100000000001",b"000100101000000001",
        -- Row: 2
        b"000000001000000010",b"000000010000000010",b"000000011000000010",b"000000100000000010",
        b"000000101000000010",b"000000110000000010",b"000001000000000010",b"000001001000000010",
        b"000001010000000010",b"000001011000000010",b"000001100000000010",b"000001110000000010",
        b"000001111000000010",b"000010000000000010",b"000010001000000010",b"000010010000000010",
        b"000010011000000010",b"000010100000000010",b"000010101000000010",b"000010110000000010",
        b"000010111000000010",b"000011000000000010",b"000011001000000010",b"000011010000000010",
        b"000011101000000010",b"000011110000000010",b"000011111000000010",b"000100000000000010",
        b"000100010000000010",b"000100011000000010",b"000100100000000010",b"000100101000000010",
        b"000100110000000010",
        -- Row: 3
        b"000000001000000011",b"000000010000000011",b"000000011000000011",b"000000100000000011",
        b"000000101000000011",b"000000110000000011",b"000000111000000011",b"000001000000000011",
        b"000001001000000011",b"000001010000000011",b"000001011000000011",b"000001100000000011",
        b"000001111000000011",b"000010000000000011",b"000010001000000011",b"000010011000000011",
        b"000010100000000011",b"000010101000000011",b"000010110000000011",b"000010111000000011",
        b"000011000000000011",b"000011101000000011",b"000011110000000011",b"000011111000000011",
        b"000100010000000011",b"000100011000000011",b"000100100000000011",b"000100101000000011",
        b"000100110000000011",
        -- Row: 4
        b"000000110000000100",b"000000111000000100",b"000001000000000100",b"000001001000000100",
        b"000001011000000100",b"000001100000000100",b"000001111000000100",b"000010000000000100",
        b"000010001000000100",b"000010011000000100",b"000010100000000100",b"000010101000000100",
        b"000011111000000100",b"000100010000000100",b"000100011000000100",b"000100100000000100",
        b"000100110000000100",
        -- Row: 5
        b"000000101000000101",b"000000110000000101",b"000000111000000101",b"000001000000000101",
        b"000001011000000101",b"000001100000000101",b"000001101000000101",b"000001111000000101",
        b"000010000000000101",b"000010100000000101",b"000010101000000101",b"000011000000000101",
        b"000011001000000101",b"000011010000000101",b"000011111000000101",b"000100000000000101",
        b"000100010000000101",b"000100011000000101",b"000100110000000101",
        -- Row: 6
        b"000000001000000110",b"000000010000000110",b"000000011000000110",b"000000100000000110",
        b"000000101000000110",b"000000110000000110",b"000001000000000110",b"000001010000000110",
        b"000001011000000110",b"000001100000000110",b"000001110000000110",b"000001111000000110",
        b"000010000000000110",b"000010010000000110",b"000010011000000110",b"000010100000000110",
        b"000010101000000110",b"000010111000000110",b"000011000000000110",b"000011001000000110",
        b"000011010000000110",b"000011110000000110",b"000011111000000110",b"000100000000000110",
        b"000100010000000110",b"000100011000000110",b"000100110000000110",
        -- Row: 7
        b"000000001000000111",b"000000010000000111",b"000000011000000111",b"000000100000000111",
        b"000000101000000111",b"000000110000000111",b"000000111000000111",b"000001000000000111",
        b"000001010000000111",b"000001011000000111",b"000001100000000111",b"000001101000000111",
        b"000001110000000111",b"000001111000000111",b"000010000000000111",b"000010010000000111",
        b"000010011000000111",b"000010100000000111",b"000010101000000111",b"000010111000000111",
        b"000011000000000111",b"000011011000000111",b"000011100000000111",b"000011101000000111",
        b"000011110000000111",b"000011111000000111",b"000100011000000111",b"000100100000000111",
        b"000100101000000111",b"000100110000000111",
        -- Row: 8
        b"000000011000001000",b"000000100000001000",b"000000101000001000",b"000001011000001000",
        b"000001110000001000",b"000001111000001000",b"000010010000001000",b"000010100000001000",
        b"000010101000001000",b"000010111000001000",b"000011000000001000",b"000011110000001000",
        b"000011111000001000",b"000100010000001000",b"000100011000001000",b"000100110000001000",
        -- Row: 9
        b"000000100000001001",b"000000101000001001",b"000000110000001001",b"000001000000001001",
        b"000001010000001001",b"000001011000001001",b"000001100000001001",b"000001101000001001",
        b"000001110000001001",b"000001111000001001",b"000010100000001001",b"000010101000001001",
        b"000010110000001001",b"000010111000001001",b"000011000000001001",b"000011111000001001",
        b"000100000000001001",b"000100011000001001",b"000100110000001001",
        -- Row: 10
        b"000000011000001010",b"000000100000001010",b"000000101000001010",b"000000110000001010",
        b"000000111000001010",b"000001000000001010",b"000001001000001010",b"000001010000001010",
        b"000001011000001010",b"000001100000001010",b"000010101000001010",b"000010110000001010",
        b"000010111000001010",b"000011000000001010",b"000011001000001010",b"000011101000001010",
        b"000011110000001010",b"000011111000001010",b"000100000000001010",b"000100011000001010",
        b"000100100000001010",
        -- Row: 11
        b"000000001000001011",b"000000010000001011",b"000000011000001011",b"000000100000001011",
        b"000001001000001011",b"000001010000001011",b"000001011000001011",b"000001100000001011",
        b"000001110000001011",b"000010000000001011",b"000010001000001011",b"000010100000001011",
        b"000010101000001011",b"000010110000001011",b"000010111000001011",b"000011000000001011",
        b"000011001000001011",b"000011010000001011",b"000011011000001011",b"000011110000001011",
        b"000011111000001011",b"000100000000001011",b"000100010000001011",b"000100011000001011",
        b"000100100000001011",
        -- Row: 12
        b"000000001000001100",b"000000010000001100",b"000000011000001100",b"000000100000001100",
        b"000000101000001100",b"000000110000001100",b"000000111000001100",b"000001000000001100",
        b"000001001000001100",b"000001010000001100",b"000001011000001100",b"000001100000001100",
        b"000001110000001100",b"000001111000001100",b"000010000000001100",b"000010001000001100",
        b"000010010000001100",b"000010011000001100",b"000010100000001100",b"000010101000001100",
        b"000010110000001100",b"000011000000001100",b"000011001000001100",b"000011010000001100",
        b"000011110000001100",b"000011111000001100",b"000100000000001100",b"000100011000001100",
        b"000100100000001100",b"000100101000001100",
        -- Row: 13
        b"000000001000001101",b"000000100000001101",b"000000101000001101",b"000001001000001101",
        b"000001011000001101",b"000001100000001101",b"000001111000001101",b"000010000000001101",
        b"000010011000001101",b"000010100000001101",b"000010101000001101",b"000010111000001101",
        b"000011000000001101",b"000011110000001101",b"000011111000001101",b"000100000000001101",
        b"000100100000001101",
        -- Row: 14
        b"000000001000001110",b"000000011000001110",b"000000100000001110",b"000000101000001110",
        b"000001000000001110",b"000001001000001110",b"000001011000001110",b"000001100000001110",
        b"000001110000001110",b"000001111000001110",b"000010000000001110",b"000010101000001110",
        b"000010110000001110",b"000010111000001110",b"000011000000001110",b"000011010000001110",
        b"000011011000001110",b"000011100000001110",b"000011101000001110",b"000011110000001110",
        b"000011111000001110",b"000100000000001110",b"000100001000001110",b"000100100000001110",
        b"000100110000001110",
        -- Row: 15
        b"000000001000001111",b"000000100000001111",b"000000101000001111",b"000000110000001111",
        b"000000111000001111",b"000001000000001111",b"000001001000001111",b"000001010000001111",
        b"000001011000001111",b"000001100000001111",b"000001101000001111",b"000001110000001111",
        b"000001111000001111",b"000010101000001111",b"000010110000001111",b"000010111000001111",
        b"000011000000001111",b"000011100000001111",b"000011101000001111",b"000011110000001111",
        b"000011111000001111",b"000100001000001111",b"000100010000001111",b"000100011000001111",
        b"000100100000001111",b"000100101000001111",b"000100110000001111",
        -- Row: 16
        b"000000001000010000",b"000000010000010000",b"000000100000010000",b"000000101000010000",
        b"000000110000010000",b"000000111000010000",b"000001000000010000",b"000001100000010000",
        b"000001101000010000",b"000001110000010000",b"000001111000010000",b"000010000000010000",
        b"000010001000010000",b"000010010000010000",b"000010101000010000",b"000010110000010000",
        b"000010111000010000",b"000011000000010000",b"000011001000010000",b"000011111000010000",
        b"000100000000010000",b"000100001000010000",b"000100010000010000",b"000100011000010000",
        -- Row: 17
        b"000000001000010001",b"000000100000010001",b"000000111000010001",b"000001000000010001",
        b"000001011000010001",b"000001101000010001",b"000001110000010001",b"000010010000010001",
        b"000010110000010001",b"000010111000010001",b"000011001000010001",b"000100000000010001",
        b"000100001000010001",
        -- Row: 18
        b"000000001000010010",b"000000010000010010",b"000000011000010010",b"000000100000010010",
        b"000000111000010010",b"000001000000010010",b"000001011000010010",b"000010000000010010",
        b"000010001000010010",b"000010010000010010",b"000010011000010010",b"000010100000010010",
        b"000010101000010010",b"000010110000010010",b"000011001000010010",b"000011100000010010",
        b"000011101000010010",b"000011110000010010",b"000011111000010010",b"000100000000010010",
        b"000100001000010010",b"000100011000010010",b"000100100000010010",b"000100101000010010",
        b"000100110000010010",
        -- Row: 19
        b"000000001000010011",b"000000111000010011",b"000001000000010011",b"000001001000010011",
        b"000001010000010011",b"000001011000010011",b"000001100000010011",b"000010010000010011",
        b"000010011000010011",b"000010100000010011",b"000010101000010011",b"000010110000010011",
        b"000010111000010011",b"000011001000010011",b"000011110000010011",b"000011111000010011",
        b"000100000000010011",b"000100001000010011",b"000100010000010011",b"000100011000010011",
        b"000100100000010011",b"000100101000010011",b"000100110000010011",
        -- Row: 20
        b"000000001000010100",b"000000010000010100",b"000000011000010100",b"000000100000010100",
        b"000000101000010100",b"000000110000010100",b"000000111000010100",b"000001000000010100",
        b"000001001000010100",b"000001010000010100",b"000001011000010100",b"000001100000010100",
        b"000001110000010100",b"000010010000010100",b"000010110000010100",b"000010111000010100",
        b"000011011000010100",b"000100000000010100",b"000100001000010100",b"000100010000010100",
        b"000100011000010100",b"000100100000010100",b"000100110000010100",
        -- Row: 21
        b"000000001000010101",b"000000010000010101",b"000000011000010101",b"000000100000010101",
        b"000000101000010101",b"000000110000010101",b"000000111000010101",b"000001010000010101",
        b"000001011000010101",b"000001100000010101",b"000001110000010101",b"000001111000010101",
        b"000010000000010101",b"000010001000010101",b"000010010000010101",b"000011011000010101",
        b"000011100000010101",b"000100000000010101",b"000100001000010101",b"000100100000010101",
        -- Row: 22
        b"000000100000010110",b"000000101000010110",b"000000110000010110",b"000001010000010110",
        b"000001011000010110",b"000001100000010110",b"000001111000010110",b"000010101000010110",
        b"000010110000010110",b"000010111000010110",b"000011000000010110",b"000011001000010110",
        b"000011011000010110",b"000011100000010110",b"000011110000010110",b"000011111000010110",
        b"000100000000010110",b"000100001000010110",b"000100100000010110",b"000100110000010110",
        -- Row: 23
        b"000000101000010111",b"000000110000010111",b"000001001000010111",b"000001010000010111",
        b"000001011000010111",b"000001100000010111",b"000001111000010111",b"000010101000010111",
        b"000010111000010111",b"000011000000010111",b"000011011000010111",b"000011110000010111",
        b"000011111000010111",b"000100000000010111",b"000100001000010111",b"000100011000010111",
        b"000100100000010111",b"000100101000010111",b"000100110000010111",
        -- Row: 24
        b"000000001000011000",b"000000010000011000",b"000000101000011000",b"000000110000011000",
        b"000001010000011000",b"000001011000011000",b"000001100000011000",b"000001110000011000",
        b"000001111000011000",b"000010000000011000",b"000010001000011000",b"000010010000011000",
        b"000010011000011000",b"000010101000011000",b"000010110000011000",b"000010111000011000",
        b"000011000000011000",b"000011001000011000",b"000011011000011000",b"000011101000011000",
        b"000011110000011000",b"000011111000011000",b"000100001000011000",b"000100011000011000",
        b"000100100000011000",b"000100110000011000",
        -- Row: 25
        b"000000001000011001",b"000000010000011001",b"000000011000011001",b"000000101000011001",
        b"000000110000011001",b"000000111000011001",b"000001010000011001",b"000001100000011001",
        b"000001111000011001",b"000010101000011001",b"000010110000011001",b"000010111000011001",
        b"000011000000011001",b"000011001000011001",b"000011010000011001",b"000011011000011001",
        b"000011100000011001",b"000011101000011001",b"000011110000011001",b"000011111000011001",
        b"000100000000011001",b"000100001000011001",b"000100011000011001",b"000100100000011001",
        b"000100101000011001",b"000100110000011001",
        -- Row: 26
        b"000000001000011010",b"000000010000011010",b"000000011000011010",b"000000100000011010",
        b"000000101000011010",b"000000110000011010",b"000000111000011010",b"000001001000011010",
        b"000001010000011010",b"000001011000011010",b"000001100000011010",b"000001101000011010",
        b"000001110000011010",b"000001111000011010",b"000010000000011010",b"000010001000011010",
        b"000010010000011010",b"000010011000011010",b"000010100000011010",b"000010101000011010",
        b"000010110000011010",b"000010111000011010",b"000011000000011010",b"000011011000011010",
        b"000011100000011010",b"000011101000011010",b"000100000000011010",b"000100001000011010",
        b"000100011000011010",b"000100100000011010",
        -- Row: 27
        b"000000001000011011",b"000000010000011011",b"000000011000011011",b"000000100000011011",
        b"000000101000011011",b"000000111000011011",b"000001000000011011",b"000001001000011011",
        b"000001010000011011",b"000001011000011011",b"000001101000011011",b"000001110000011011",
        b"000001111000011011",b"000010000000011011",b"000010001000011011",b"000010010000011011",
        b"000010011000011011",b"000010100000011011",b"000010101000011011",b"000010110000011011",
        b"000010111000011011",b"000011010000011011",b"000011011000011011",b"000011100000011011",
        b"000011101000011011",b"000011110000011011",b"000100001000011011",b"000100010000011011",
        b"000100100000011011",b"000100101000011011",
        -- Row: 28
        b"000000011000011100",b"000000100000011100",b"000001000000011100",b"000001001000011100",
        b"000001010000011100",b"000001110000011100",b"000001111000011100",b"000010000000011100",
        b"000010010000011100",b"000010011000011100",b"000010101000011100",b"000010110000011100",
        b"000011011000011100",b"000011100000011100",b"000100100000011100",b"000100101000011100",
        b"000100110000011100"
        -- Row: 29
	        );
	
    signal track_1_free_pos_mem : track_1_free_pos_mem_t := track_1_free_pos_mem_c;
    signal track_2_free_pos_mem : track_2_free_pos_mem_t := track_2_free_pos_mem_c;
    signal track_3_free_pos_mem : track_3_free_pos_mem_t := track_3_free_pos_mem_c;
    signal track_4_free_pos_mem : track_4_free_pos_mem_t := track_4_free_pos_mem_c;

begin 
    
    --****************************
    --* Random number generation *
    --****************************
    free_pos_lmt <= 
    to_signed(913,11)   when (NEXT_TRACK(1 downto 0) = "00") else
    to_signed(886,11)   when (NEXT_TRACK(1 downto 0) = "01") else
    to_signed(932,11)   when (NEXT_TRACK(1 downto 0) = "10") else
    to_signed(660,11)   when (NEXT_TRACK(1 downto 0) = "11") else
    (others => '0');
    
    -- Counter to take bits from
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                free_pos_cnt <= (others => '0');
            elsif (free_pos_cnt >= free_pos_lmt) then
                free_pos_cnt <= (others => '0');
            else
                free_pos_cnt <= free_pos_cnt + 1;
            end if;
        end if;
    end process;
    
    --*********************************************************
    --* RND_GOAL_POS : Random, free position in current track *
    --*********************************************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                RND_GOAL_POS <= track_1_free_pos_mem(0);
            else
                case sel_track is
                    when "00" =>
                        RND_GOAL_POS <= track_1_free_pos_mem(to_integer(free_pos_cnt));
                    when "01" =>
                        RND_GOAL_POS <= track_2_free_pos_mem(to_integer(free_pos_cnt));
                    when "10" =>
                        RND_GOAL_POS <= track_3_free_pos_mem(to_integer(free_pos_cnt));
                    when "11" =>
                        RND_GOAL_POS <= track_4_free_pos_mem(to_integer(free_pos_cnt));
                    when others =>
                        RND_GOAL_POS <= track_4_free_pos_mem(to_integer(free_pos_cnt));
                        --null;
                end case;
            end if;
        end if;
    end process;
    
	--*****************************
    --* IR : Instruction Register *
    --*****************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                IR <= (others => '0');
            elsif (FB = "001") then
                IR <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;
    
    OP <= IR(17 downto 13);   -- Operation    
    GRX <= IR(12 downto 10);  -- Register    
    M <= IR(9 downto 8);      -- Addressing mode        
    ADDR <= IR(7 downto 0);   -- Address field

    -- FB = "010" UNUSED (CAN'T WRITE TO PM)
    
    --************************
    --* PC : Program Counter *
    --************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                PC <= (others => '0');
            elsif (FB = "011") then
                PC <= DATA_BUS(7 downto 0);
            elsif (P = '1') then
                PC <= PC + 1;
            else
                null;
            end if;
        end if;
    end process;

    --*********************************************
    --* WON : Signal for when goal pos was found. *
    --*********************************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                WON <= '0';
            elsif (FB = "100") then
                WON <= DATA_BUS(0);
            else
                null;
            end if;
        end if;
    end process; 

    --*********************************
    --* SCORE : Current player score. *
    --*********************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                SCORE <= (others => '0');
            elsif (FB = "101") then
                SCORE <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process; 
    
    --****************************
    --* GR0 : General Register 0 *
    --****************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                GR0 <= (others => '0');
            elsif (S = '1') then
                if (M = "00") then
                    GR0 <= DATA_BUS;
                else 
                    null;
                end if;
            elsif (FB = "110" and GRX = "000") then
                GR0 <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;
    
    --****************************
    --* GR1 : General Register 1 *
    --****************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                GR1 <= (others => '0');
            elsif (S = '1') then
                if (M = "01") then
                    GR1 <= DATA_BUS;
                else 
                    null;
                end if;
            elsif (FB = "110" and GRX = "001") then
                GR1 <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;
    
    --****************************
    --* GR2 : General Register 2 *
    --****************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                GR2 <= (others => '0');
            elsif (S = '1') then
                if (M = "10") then
                    GR2 <= DATA_BUS;
                else 
                    null;
                end if;
            elsif (FB = "110" and GRX = "010") then
                GR2 <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;
    
    --****************************
    --* GR3 : General Register 3 *
    --****************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                GR3 <= (others => '0');
            elsif (S = '1') then
                if (M = "11") then
                    GR3 <= DATA_BUS;
                else 
                    null;
                end if;
            elsif (FB = "110" and GRX = "011") then
                GR3 <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;
    
    --************************************
    --* GOAL_POS : Goal Position Register *
    --************************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                GOAL_POS <= (others => '0');
            elsif (FB = "110" and GRX = "100") then
                GOAL_POS <= DATA_BUS;
            else
                null;
            end if;
        end if;
    end process;


    ----*****************************************
    ----* NEXT_TRACK : Track-selection Register *
    ----*****************************************  
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                SEL_TRACK <= "00";
                NEXT_TRACK <= (others => '1');
                dly_cnt <= to_unsigned(0,3);
            -- In process of changing track, locking keyboard.
            elsif (dly_cnt = "000" and FB = "110" and GRX = "101") then
                NEXT_TRACK <= DATA_BUS; 
                dly_cnt <= to_unsigned(1,3);
            elsif (dly_cnt = "001") then
                dly_cnt <= to_unsigned(2,3);
            elsif (dly_cnt = "010") then
                dly_cnt <= to_unsigned(3,3);
            -- Changing track and requesting updated sound icon (in key pressed section).
            elsif (dly_cnt = "011") then
                dly_cnt <= to_unsigned(4,3);
                SEL_TRACK <= NEXT_TRACK(1 downto 0);
            elsif (dly_cnt = "100") then
                dly_cnt <= to_unsigned(5,3);
            elsif (dly_cnt = "101") then
                dly_cnt <= to_unsigned(0,3);            
            else
                null;
            end if;
        end if;
    end process;    

    --FB = "110" & GRX = "110" UNUSED
    --FB = "110" & GRX = "111" UNUSED
    
    --*****************************************
    --* ASR : Program Memory Address Register *
    --*****************************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                ASR <= (others => '0');
            elsif (FB = "111") then 
                ASR <= DATA_BUS(7 downto 0);
            end if;
        end if;
    end process;
   
   
    --*******************************
    --* uPC : Micro Program Counter *
    --*******************************
    process(clk)
    begin
    if rising_edge(clk) then
        if (rst = '1') then
            uPC <= (others => '0');
        else
            case SEQ is
                when "0000" =>
                    uPC <= uPC + 1;
                when "0001" => 
                    uPC <= uAddr_instr(to_integer(unsigned(OP)));
                when "0010" =>
                    case M is
                        when "00" =>
                            uPC <= "0000011"; -- "Direct adressering" uAddr
                        when "01" => 
                            uPC <= "0000100"; -- "Immediate operand" uAddr
                        when "10" => 
                            uPC <= "0000101"; -- "Indirect adressering" uAddr
                        when "11" => 
                            uPC <= "0000111"; -- "Indexed adressering" uAddr
                        when others => 
                            uPC <= (others => '0');
                    end case;
                when "0011" =>
                    uPC <= (others => '0');
                when "0100" =>
                    if (flag_Z = '0') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if;        
                when "0101" =>          
                    uPC <= MICROADDR;
                when "0110" =>
                    if (flag_S = '0') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if; 
                -- "0111" UNUSED (Subroutine-related)
                when "1000" =>
                    if (flag_Z = '1') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                   end if;
                when "1001" =>
                    if (flag_N = '1') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if;
                --when "1010" =>
                --    if (flag_C = '1') then
                --        uPC <= MICROADDR;
                --    else 
                --        uPC <= uPC + 1;
                --    end if;
                when "1011" =>
                    if (flag_O = '1') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if;
                when "1100" =>
                    if (flag_L = '1') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if;  
                when "1101" =>  -- Used in BCT (branch on continue).
                    if (flag_G = '1') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if; 
                when "1110" =>
                    if (flag_O = '0') then
                        uPC <= MICROADDR;
                    else 
                        uPC <= uPC + 1;
                    end if;  
               --when "1111" => ***UNUSED***
               --     uPC <= (others => '0'); -- SHOULD ALSO HALT EXECUTION   
               when others =>
                    null;
            end case; 
        end if;
    end if;
    end process;
    
    --******************************
    --* Goal position reached flag *
    --******************************
    flag_G <= '1' when (CURR_POS = GOAL_POS) else '0';  
    
    --*****************************
    --* Showing goal message flag *
    --*****************************
    flag_S <= '1' when (showing_goal_msg = '1') else '0';  
    
    --*******************************
    --* ALU : Arithmetic Logic Unit *
    --*******************************
    process(clk)
    begin
    if rising_edge(clk) then
        if rst = '1' then
            AR <= (others => '0');
            --flag_C <= '0';
            --flag_O <= '0';
        else
            case ALU is
                when "0000" =>  -- NO FUNCTION (No flags) 
                    null;      
                when "0001" => -- AR := DATA_BUS (No flags)
                    AR <= DATA_BUS;      
                --when "0010" =>  -- ONES' COMPLEMENT, (No flags) ***UNUSED***
                when "0011" =>  -- SET TO ZERO (Z/N)            ***UNUSED***
                    AR <= (others => '0');   
                when "0100" => -- AR := AR + DATA_BUS (Z/N/O/C)
                    AR <= AR + DATA_BUS;
                    -- SHOULD SET OVERFLOW AND CARRY AS WELL   
                when "0101" => -- AR := AR - DATA_BUS (Z/N/O/C)
                    AR <= AR - DATA_BUS;
                    -- SHOULD SET OVERFLOW AND CARRY AS WELL       
                when "0110" => -- AR := AR and DATA_BUS (Z/N)
                    AR <= AR and DATA_BUS;        
                 --when "0111" => -- AR := AR or DATA_BUS (Z/N)       ***UNUSED***
                 --   AR <= AR or DATA_BUS;     
                when "1000" => -- AR := 1 (Z/N)
                    AR <= to_signed(1,18);                      
                --when "1001" => -- AR LSL, zero is shifted in, bit shifted out to C. (Z/N(C) ***UNUSED***
                --    AR <= AR(16 downto 0) & '0';
                --    flag_C <= AR(17);   
                --when "1010" => -- AR LSL, 32-bit,                   ***UNUSED*** 
                --when "1011" => -- AR ASR, sign bit is shifted in, bit shifted out to C. (Z/N/C) ***UNUSED***
                --    AR <= AR(17) & AR(17 downto 1);
                --    flag_C <= AR(0);
                --when "1100" => -- ARHR ASR,                         ***UNUSED***
                when "1101" => -- AR LSR, zero is shifted in, bit shifted out to C. (Z/N/C)
                    AR <= '0' & AR(17 downto 1);
                    --flag_C <= AR(0);
                --when "1110" => -- Rotate AR to the left,            ***UNUSED***
                --when "1111" => -- Rotate ARHR to the left (32-bit), ***UNUSED***
                when others =>
                    null;
     
            end case;
        end if;
    end if;
    end process;
    flag_Z <= '1' when (AR = to_signed(0,18)) else '0';
    flag_N <= '1' when (AR < to_signed(0,18)) else '0';
    flag_C <= '0'; -- NOT BEING DETECTED ATM, MIGHT HAVE TO IMPLEMENT INSIDE ALU PROCESS
    flag_O <= '0'; -- NOT BEING DETECTED ATM, MIGHT HAVE TO IMPLEMENT INSIDE ALU PROCESS

    --*********************
    --* LC : Loop Counter *
    --*********************
    process(clk)
    begin
    if rising_edge(clk) then
        if rst = '1' then
            LC_cnt <= (others => '0');
        else
            if (LC = "01" and LC_cnt > 0) then
                LC_cnt <= LC_cnt - 1;
            elsif (LC = "10") then
                LC_cnt <= to_signed(0,9) & DATA_BUS(7 downto 0);
            elsif (LC = "11") then
                LC_cnt <= to_signed(0,10) & signed(MICROADDR);
            else
                null;
            end if;
        end if;
    end if;
    end process;
    
    flag_L <= '1' when (LC_cnt = 0) else '0';

    --***********************
    --* Data Bus Assignment *
    --***********************
    DATA_BUS <= 
    to_signed(0,10) & IR(7 downto 0)    when (TB = "001") else  -- ADR
    PM                                  when (TB = "010") else
    to_signed(0,10) & PC                when (TB = "011") else
    AR                                  when (TB = "100") else
    SCORE                               when (TB = "101") else
    GR0                                 when (TB = "110" and GRX = "000") else 
    GR1                                 when (TB = "110" and GRX = "001") else 
    GR2                                 when (TB = "110" and GRX = "010") else 
    GR3                                 when (TB = "110" and GRX = "011") else
    RND_GOAL_POS                        when (TB = "110" and GRX = "100") else
    NEXT_TRACK                          when (TB = "110" and GRX = "101") else 
    --NULL                                when (TB = "110" and GRX = "110") else 
    --NULL                                when (TB = "110" and GRX = "111") else 
    to_signed(0,16) & SEL_TRACK         when (TB = "110" and GRX = "111") else
    to_signed(0,10) & ASR               when (TB = "111") else
    DATA_BUS;
    
    --*************************
    --* PS2cmd Interpretation *
    --*************************
    process(clk)
    begin
        if rising_edge(clk) then
            if (rst = '1') then
                CURR_POS <= "000000001000000001";
                NEXT_POS <= "000000001000000001";
                MOVE_REQ <= '0';
                UPD_SOUND_ICON <= '0';
                DISP_GOAL_POS <= '0';
                SEL_SOUND <= '0';
            else
                if (move_resp = '1') then
                    CURR_POS <= NEXT_POS;
                end if;
                UPD_SOUND_ICON <= '0';
                MOVE_REQ <= '0';
                -- We're changing track, send move_req back to start.
                if (dly_cnt = 0 and FB = "110" and GRX = "101") then  
                    NEXT_POS <= "000000001000000001";
                    MOVE_REQ <= '1';
                -- Not in locked mode, check for key pressed.
                elsif (dly_cnt = 0) then
                    case key_code is
                        when "001" =>  -- UP (W)
                            NEXT_XPOS <= CURR_XPOS;
                            NEXT_YPOS <= CURR_YPOS - 1;
                            MOVE_REQ <= '1';
                        when "010" =>  -- LEFT (A)
                            NEXT_YPOS <= CURR_YPOS;
                            NEXT_XPOS <= CURR_XPOS - 1;
                            MOVE_REQ <= '1';
                        when "011" =>  -- DOWN (S)
                            NEXT_XPOS <= CURR_XPOS;
                            NEXT_YPOS <= CURR_YPOS + 1;
                            MOVE_REQ <= '1';
                        when "100" =>  -- RIGHT (D)
                            NEXT_YPOS <= CURR_YPOS;
                            NEXT_XPOS <= CURR_XPOS + 1;
                            MOVE_REQ <= '1';
                        when "101" => -- DISPLAY GOAL POS TOGGLE (G)
                            DISP_GOAL_POS <= not DISP_GOAL_POS;
                        when "110" => -- SOUND TOGGLE (SPACE)
                            SEL_SOUND <= not SEL_SOUND;
                            UPD_SOUND_ICON <= '1';
                        when others =>
                            null;
                    end case;
                -- In locked mode, don't check for key pressed.
                -- Time to update sound icon
                elsif (dly_cnt = 3) then
                    UPD_SOUND_ICON <= '1';
                -- Do nothing, GPU busy
                else    
                    null;
                end if;
            end if;
        end if;
    end process;
 
    --*******************************
    --* Outgoing signals assignment *
    --*******************************
    pAddr <= ASR when (ASR >= to_signed(0,8) and ASR <= to_signed(13,8)) else to_signed(0,8);
    uAddr <= uPC; 
    curr_pos_out <= CURR_POS;
    next_pos_out <= NEXT_POS;
    goal_pos_out <= GOAL_POS;
    sel_track_out <= unsigned(SEL_TRACK);
    sel_sound_out <= SEL_SOUND;
    move_req_out <= MOVE_REQ;
    upd_sound_icon_out <= UPD_SOUND_ICON;
    goal_reached_out <= WON;
    disp_goal_pos_out <= DISP_GOAL_POS;
    score_out <= unsigned(SCORE(5 downto 0));

end Behavioral;


