--------------------------------------------------------------------------------
-- PIC MEM
-- ZigSound
-- 04-apr-2017
-- Version 0.1


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity PIC_MEM is
	port(
        clk		        	: in std_logic;
        rst		            : in std_logic;
        -- CPU
        sel_track       	: in unsigned(1 downto 0);
        -- GPU
        we		        	: in std_logic;
        data_nextpos    	: out unsigned(7 downto 0);
        addr_nextpos    	: in unsigned(10 downto 0);
        data_change	    	: in unsigned(7 downto 0);
        addr_change	    	: in unsigned(10 downto 0);
        -- VGA MOTOR
        data_vga        	: out unsigned(7 downto 0);
        addr_vga	    	: in unsigned(10 downto 0)
	);

end PIC_MEM;
	
-- Architecture
architecture Behavioral of PIC_MEM is

    -- Track memory type
    type ram_t is array (0 to 1199) of unsigned(7 downto 0);
    -- Maximum array length is 2048, change when adding/deleting from ram_t.

    -- TRACK 1 initialization
    signal track_1 : ram_t := (
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 0
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 0
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 0
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 0
        x"18",x"1F",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 1
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 1
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 1
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 1
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 2
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 2
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 2
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 2
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 3
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 3
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 3
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 3
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 4
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 4
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 4
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 4
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 5
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 5
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 5
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 5
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 6
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 6
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 6
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 6
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 7
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 7
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 7
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 7
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 8
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 8
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 8
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 8
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 9
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 9
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 9
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 9
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 10
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 10
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 10
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 10
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 11
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 11
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 11
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 11
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 12
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 12
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 12
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 12
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 13
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 13
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 13
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 13
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 14
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 14
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 14
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 14
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 15
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 15
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 15
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 15
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 16
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 16
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 16
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 16
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 17
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 17
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 17
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 17
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 18
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 18
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 18
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 18
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 19
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 19
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 19
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 19
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 20
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 20
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 20
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 20
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 21
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 21
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 21
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 21
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 22
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 22
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 22
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 22
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 23
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 23
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 23
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 23
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 24
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 24
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 24
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 24
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 25
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 25
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 25
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 25
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 26
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 26
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 26
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 26
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 27
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 27
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 27
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 27
        x"18",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 28
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 28
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- Row 28
        x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"18", -- Row 28
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 29
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 29
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18", -- Row 29
        x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18",x"18"  -- Row 29
        );
        
    -- TRACK 2 initialization
    signal track_2 : ram_t := (0 => x"1F", others => (others => '0')); 
    
    -- TRACK 3 initialization
    signal track_3 : ram_t := (0 => x"1F", others => (others => '0')); 


begin

    -- Checks if write enable, in that case makes changes to memory using 
    -- addr_change and data_change.
    process(clk)
    begin
    if rising_edge(clk) then
        if (rst = '1') then
            null;
        elsif (we = '1') then
            track_1(1) <= x"02";
            case sel_track is
                when "01" =>
                    track_1(to_integer(addr_change)) <= data_change;
                when "10" =>
                    track_2(to_integer(addr_change)) <= data_change;
                when "11" =>
                    track_3(to_integer(addr_change)) <= data_change;
                when others =>
                    null;
            end case;
        else
            track_1(0) <= x"01";
        end if;  
    end if;
    end process;

    -- Sets data_nextpos to data at addr_nextpos and data_vga to data at addr_vga.
    with sel_track select
        data_nextpos <= 
        track_1(to_integer(addr_nextpos)) when "01",
        track_2(to_integer(addr_nextpos)) when "10",
        track_3(to_integer(addr_nextpos)) when "11",
        "00000000" when others;
    with sel_track select
        data_vga <= 
        track_1(to_integer(addr_vga)) when "01",
        track_2(to_integer(addr_vga)) when "10",
        track_3(to_integer(addr_vga)) when "11",
        "00000000" when others;

end Behavioral;

