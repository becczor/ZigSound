--------------------------------------------------------------------------------
-- PIC MEM
-- ZigSound
-- 04-apr-2017
-- Version 0.1


-- library declaration
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;            -- basic IEEE library
use IEEE.NUMERIC_STD.ALL;               -- IEEE library for the unsigned type


-- entity
entity PIC_MEM is
	port(
        clk		        	: in std_logic;
        rst		            : in std_logic;
        -- CPU
        sel_track       	: in unsigned(1 downto 0);
        -- GPU
        we		        	: in std_logic;
        data_nextpos    	: out unsigned(7 downto 0);
        addr_nextpos    	: in unsigned(10 downto 0);
        data_change	    	: in unsigned(7 downto 0);
        addr_change	    	: in unsigned(10 downto 0);
        -- VGA MOTOR
        data_vga        	: out unsigned(7 downto 0);
        addr_vga	    	: in unsigned(10 downto 0)
	);

end PIC_MEM;
	
-- Architecture
architecture Behavioral of PIC_MEM is


    -- Track memory type
    type ram_t is array (0 to 4799) of unsigned(7 downto 0);
    -- Track initialization
    signal track : ram_t := (
        --***********
        --* TRACK 1 *
        --***********
        x"06",x"06",x"06",x"07",x"06",x"06",x"07",x"07",x"07",x"06",x"06",x"07",x"06",x"06",x"07",x"06",x"06",x"06",x"06",x"07",x"07",x"06",x"06",x"07",x"07",x"07",x"06",x"06",x"06",x"06",x"07",x"06",x"07",x"06",x"06",x"06",x"06",x"06",x"06",x"06",
        x"07",x"03",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"07",
        x"06",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"07",x"06",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
        x"07",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"06",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"06",
        x"07",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"06",
        x"07",x"07",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"06",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"00",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"06",
        x"07",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"07",x"00",x"00",x"06",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"07",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"07",x"00",x"07",
        x"07",x"00",x"00",x"00",x"06",x"00",x"06",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"07",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"06",x"07",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"06",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"07",
        x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"06",x"06",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"07",x"00",x"07",
        x"06",x"00",x"00",x"00",x"07",x"06",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"06",
        x"07",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",
        x"06",x"00",x"07",x"06",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"04",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"07",x"00",x"00",x"07",
        x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"07",
        x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"06",
        x"06",x"00",x"00",x"00",x"00",x"06",x"07",x"00",x"00",x"00",x"06",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"07",x"06",
        x"06",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"06",x"00",x"00",x"06",x"00",x"00",x"00",x"06",x"00",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"07",x"00",x"00",x"00",x"00",x"00",x"07",x"06",
        x"06",x"06",x"07",x"07",x"06",x"06",x"06",x"07",x"06",x"06",x"07",x"07",x"06",x"06",x"07",x"06",x"06",x"06",x"07",x"07",x"06",x"06",x"07",x"07",x"06",x"06",x"07",x"06",x"06",x"06",x"07",x"07",x"06",x"06",x"06",x"06",x"06",x"06",x"06",x"0C",
        --***********
        --* TRACK 2 *
        --***********
        x"09",x"08",x"08",x"09",x"09",x"08",x"08",x"08",x"09",x"09",x"08",x"08",x"09",x"08",x"08",x"08",x"09",x"09",x"08",x"08",x"08",x"09",x"09",x"09",x"08",x"08",x"09",x"08",x"08",x"08",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"09",x"08",x"08",
        x"08",x"03",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"09",x"09",
        x"08",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"08",
        x"08",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"08",
        x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"04",x"01",x"09",
        x"08",x"01",x"09",x"01",x"08",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"08",
        x"08",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"08",x"09",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",
        x"08",x"01",x"08",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"04",x"08",x"01",x"01",x"01",x"01",x"01",x"08",
        x"08",x"01",x"01",x"01",x"01",x"08",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"08",x"01",x"01",x"01",x"09",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",
        x"09",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"08",
        x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"09",
        x"08",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",
        x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"09",
        x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"08",
        x"08",x"01",x"08",x"09",x"04",x"01",x"01",x"01",x"04",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"09",x"01",x"01",x"01",x"01",x"08",
        x"09",x"01",x"01",x"01",x"08",x"01",x"01",x"08",x"09",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"08",
        x"08",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"08",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"08",x"08",x"01",x"08",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",
        x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"08",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",
        x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"08",x"01",x"01",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"08",x"08",x"01",x"01",x"01",x"01",x"01",x"08",
        x"09",x"01",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"04",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"09",
        x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"09",
        x"08",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"04",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",
        x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"09",
        x"08",x"09",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"08",
        x"09",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"08",x"01",x"04",x"01",x"01",x"01",x"08",
        x"08",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"08",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",
        x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"09",x"01",x"01",x"01",x"08",x"01",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"01",x"08",
        x"09",x"01",x"08",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"08",x"01",x"01",x"01",x"08",x"09",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"09",x"08",x"01",x"08",
        x"08",x"09",x"01",x"01",x"01",x"09",x"08",x"04",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",x"01",x"01",x"01",x"01",x"01",x"01",x"09",x"08",
        x"09",x"08",x"08",x"09",x"08",x"08",x"09",x"08",x"08",x"09",x"09",x"08",x"08",x"09",x"08",x"08",x"08",x"08",x"09",x"08",x"08",x"08",x"09",x"08",x"08",x"09",x"08",x"09",x"09",x"08",x"08",x"09",x"08",x"08",x"09",x"09",x"09",x"09",x"08",x"0C",
        --***********
        --* TRACK 3 *
        --***********
        x"0A",x"0A",x"0B",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
        x"0B",x"03",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"0B",x"05",x"0B",x"0A",
        x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",
        x"0A",x"0B",x"02",x"02",x"02",x"05",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"0B",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0A",x"02",x"02",x"02",x"05",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0A",
        x"0A",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"0A",
        x"0B",x"0A",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0B",
        x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"0A",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"0A",x"05",x"02",x"0A",x"0B",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0B",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"0B",
        x"0A",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",
        x"0A",x"0A",x"0B",x"02",x"02",x"02",x"02",x"05",x"0A",x"0A",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"05",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0B",x"0A",x"0B",x"0B",x"0B",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0C",
        --***********
        --* TRACK 4 *
        --***********
        x"0A",x"0A",x"0B",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",
        x"0B",x"03",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"0B",x"05",x"0B",x"0A",
        x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",
        x"0A",x"0B",x"02",x"02",x"02",x"05",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"0B",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0A",x"02",x"02",x"02",x"05",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0A",
        x"0A",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"0A",
        x"0B",x"0A",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0B",
        x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"0A",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"0A",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"0A",x"05",x"02",x"0A",x"0B",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"0B",x"02",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",x"02",x"0B",
        x"0A",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"0A",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"0A",
        x"0B",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"02",x"02",x"0B",
        x"0A",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0B",x"02",x"0A",
        x"0A",x"0A",x"0B",x"02",x"02",x"02",x"02",x"05",x"0A",x"0A",x"02",x"02",x"02",x"02",x"05",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"02",x"0A",x"05",x"02",x"02",x"02",x"0A",x"02",x"02",x"02",x"02",x"0A",
        x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0B",x"0A",x"0B",x"0B",x"0B",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0B",x"0B",x"0A",x"0A",x"0A",x"0B",x"0A",x"0A",x"0A",x"0A",x"0A",x"0A",x"0C"
        );
        

begin

    -- Checks if write enable, in that case makes changes to memory using 
    -- addr_change and data_change.
    process(clk)
    begin
    if rising_edge(clk) then
        if (we = '1') then
            track(to_integer(sel_track*to_unsigned(1200,11) + addr_change)) <= data_change;
        else
            null;
        end if;
        -- Uses sel_track to get correct track index to then set data out to correct tile
        data_vga <= track(to_integer(sel_track*to_unsigned(1200,11) + addr_vga));
        data_nextpos <= track(to_integer(sel_track*to_unsigned(1200,11) + addr_nextpos));
    end if;
    end process;

end Behavioral;

